library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity testbench is
end testbench ;
architecture Behavioral of testbench is
constant CLK_PERIOD : time := 2 ns; -- Clock period
signal clk_tb : std_logic := '0';
signal x_0_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_1_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_2_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_3_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_4_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_5_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_6_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_7_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_8_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_9_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_10_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_11_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_12_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_13_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_14_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_15_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_16_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_17_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_18_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_19_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_20_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_21_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_22_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_23_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_24_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_25_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_26_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_27_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_28_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_29_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_30_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_31_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_32_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_33_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_34_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_35_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_36_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_37_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_38_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_39_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_40_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_41_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_42_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_43_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_44_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_45_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_46_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_47_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_48_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_49_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_50_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_51_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_52_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_53_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_54_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_55_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_56_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_57_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_58_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_59_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_60_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_61_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_62_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_63_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_64_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_65_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_66_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_67_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_68_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_69_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_70_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_71_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_72_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_73_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_74_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_75_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_76_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_77_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_78_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_79_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_80_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_81_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_82_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_83_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_84_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_85_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_86_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_87_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_88_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_89_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_90_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_91_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_92_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_93_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_94_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_95_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_96_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_97_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_98_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_99_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_100_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_101_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_102_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_103_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_104_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_105_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_106_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_107_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_108_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_109_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_110_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_111_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_112_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_113_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_114_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_115_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_116_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_117_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_118_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_119_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_120_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_121_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_122_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_123_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_124_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_125_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_126_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_127_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_128_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_129_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_130_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_131_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_132_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_133_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_134_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_135_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_136_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_137_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_138_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_139_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_140_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_141_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_142_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_143_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_144_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_145_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_146_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_147_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_148_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_149_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_150_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_151_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_152_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_153_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_154_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_155_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_156_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_157_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_158_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_159_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_160_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_161_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_162_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_163_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_164_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_165_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_166_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_167_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_168_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_169_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_170_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_171_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_172_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_173_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_174_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_175_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_176_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_177_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_178_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_179_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_180_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_181_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_182_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_183_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_184_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_185_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_186_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_187_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_188_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_189_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_190_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_191_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_192_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_193_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_194_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_195_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_196_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_197_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_198_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_199_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_200_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_201_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_202_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_203_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_204_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_205_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_206_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_207_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_208_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_209_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_210_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_211_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_212_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_213_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_214_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_215_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_216_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_217_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_218_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_219_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_220_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_221_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_222_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_223_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_224_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_225_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_226_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_227_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_228_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_229_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_230_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_231_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_232_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_233_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_234_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_235_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_236_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_237_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_238_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_239_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_240_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_241_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_242_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_243_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_244_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_245_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_246_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_247_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_248_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_249_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_250_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_251_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_252_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_253_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_254_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_255_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_256_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_257_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_258_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_259_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_260_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_261_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_262_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_263_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_264_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_265_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_266_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_267_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_268_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_269_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_270_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_271_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_272_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_273_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_274_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_275_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_276_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_277_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_278_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_279_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_280_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_281_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_282_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_283_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_284_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_285_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_286_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_287_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_288_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_289_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_290_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_291_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_292_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_293_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_294_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_295_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_296_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_297_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_298_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_299_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_300_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_301_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_302_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_303_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_304_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_305_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_306_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_307_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_308_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_309_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_310_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_311_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_312_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_313_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_314_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_315_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_316_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_317_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_318_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_319_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_320_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_321_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_322_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_323_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_324_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_325_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_326_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_327_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_328_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_329_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_330_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_331_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_332_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_333_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_334_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_335_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_336_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_337_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_338_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_339_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_340_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_341_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_342_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_343_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_344_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_345_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_346_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_347_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_348_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_349_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_350_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_351_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_352_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_353_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_354_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_355_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_356_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_357_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_358_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_359_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_360_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_361_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_362_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_363_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_364_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_365_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_366_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_367_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_368_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_369_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_370_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_371_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_372_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_373_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_374_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_375_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_376_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_377_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_378_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_379_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_380_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_381_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_382_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_383_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_384_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_385_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_386_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_387_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_388_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_389_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_390_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_391_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_392_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_393_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_394_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_395_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_396_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_397_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_398_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_399_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_400_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_401_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_402_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_403_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_404_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_405_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_406_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_407_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_408_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_409_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_410_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_411_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_412_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_413_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_414_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_415_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_416_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_417_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_418_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_419_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_420_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_421_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_422_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_423_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_424_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_425_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_426_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_427_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_428_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_429_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_430_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_431_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_432_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_433_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_434_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_435_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_436_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_437_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_438_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_439_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_440_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_441_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_442_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_443_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_444_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_445_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_446_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_447_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_448_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_449_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_450_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_451_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_452_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_453_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_454_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_455_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_456_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_457_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_458_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_459_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_460_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_461_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_462_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_463_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_464_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_465_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_466_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_467_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_468_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_469_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_470_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_471_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_472_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_473_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_474_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_475_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_476_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_477_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_478_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_479_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_480_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_481_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_482_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_483_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_484_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_485_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_486_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_487_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_488_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_489_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_490_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_491_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_492_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_493_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_494_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_495_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_496_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_497_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_498_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_499_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_500_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_501_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_502_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_503_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_504_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_505_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_506_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_507_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_508_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_509_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_510_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_511_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_512_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_513_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_514_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_515_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_516_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_517_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_518_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_519_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_520_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_521_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_522_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_523_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_524_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_525_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_526_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_527_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_528_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_529_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_530_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_531_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_532_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_533_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_534_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_535_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_536_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_537_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_538_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_539_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_540_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_541_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_542_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_543_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_544_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_545_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_546_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_547_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_548_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_549_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_550_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_551_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_552_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_553_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_554_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_555_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_556_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_557_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_558_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_559_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_560_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_561_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_562_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_563_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_564_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_565_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_566_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_567_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_568_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_569_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_570_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_571_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_572_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_573_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_574_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_575_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_576_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_577_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_578_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_579_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_580_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_581_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_582_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_583_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_584_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_585_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_586_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_587_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_588_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_589_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_590_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_591_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_592_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_593_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_594_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_595_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_596_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_597_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_598_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_599_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_600_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_601_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_602_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_603_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_604_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_605_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_606_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_607_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_608_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_609_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_610_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_611_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_612_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_613_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_614_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_615_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_616_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_617_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_618_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_619_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_620_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_621_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_622_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_623_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_624_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_625_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_626_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_627_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_628_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_629_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_630_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_631_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_632_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_633_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_634_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_635_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_636_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_637_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_638_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_639_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_640_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_641_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_642_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_643_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_644_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_645_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_646_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_647_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_648_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_649_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_650_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_651_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_652_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_653_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_654_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_655_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_656_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_657_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_658_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_659_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_660_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_661_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_662_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_663_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_664_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_665_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_666_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_667_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_668_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_669_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_670_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_671_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_672_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_673_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_674_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_675_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_676_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_677_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_678_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_679_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_680_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_681_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_682_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_683_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_684_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_685_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_686_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_687_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_688_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_689_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_690_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_691_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_692_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_693_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_694_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_695_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_696_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_697_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_698_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_699_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_700_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_701_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_702_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_703_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_704_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_705_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_706_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_707_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_708_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_709_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_710_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_711_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_712_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_713_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_714_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_715_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_716_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_717_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_718_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_719_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_720_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_721_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_722_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_723_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_724_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_725_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_726_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_727_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_728_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_729_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_730_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_731_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_732_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_733_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_734_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_735_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_736_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_737_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_738_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_739_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_740_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_741_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_742_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_743_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_744_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_745_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_746_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_747_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_748_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_749_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_750_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_751_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_752_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_753_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_754_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_755_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_756_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_757_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_758_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_759_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_760_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_761_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_762_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_763_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_764_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_765_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_766_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_767_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_768_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_769_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_770_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_771_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_772_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_773_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_774_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_775_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_776_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_777_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_778_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_779_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_780_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_781_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_782_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal x_783_tb  : STD_LOGIC_VECTOR(15 downto 0);
signal y_tb  : STD_LOGIC_VECTOR(3 downto 0);
begin
	dut: entity work.lstm
	Port map (
clk => clk_tb ,
	x_0 => x_0_tb,
	x_1 => x_1_tb,
	x_2 => x_2_tb,
	x_3 => x_3_tb,
	x_4 => x_4_tb,
	x_5 => x_5_tb,
	x_6 => x_6_tb,
	x_7 => x_7_tb,
	x_8 => x_8_tb,
	x_9 => x_9_tb,
	x_10 => x_10_tb,
	x_11 => x_11_tb,
	x_12 => x_12_tb,
	x_13 => x_13_tb,
	x_14 => x_14_tb,
	x_15 => x_15_tb,
	x_16 => x_16_tb,
	x_17 => x_17_tb,
	x_18 => x_18_tb,
	x_19 => x_19_tb,
	x_20 => x_20_tb,
	x_21 => x_21_tb,
	x_22 => x_22_tb,
	x_23 => x_23_tb,
	x_24 => x_24_tb,
	x_25 => x_25_tb,
	x_26 => x_26_tb,
	x_27 => x_27_tb,
	x_28 => x_28_tb,
	x_29 => x_29_tb,
	x_30 => x_30_tb,
	x_31 => x_31_tb,
	x_32 => x_32_tb,
	x_33 => x_33_tb,
	x_34 => x_34_tb,
	x_35 => x_35_tb,
	x_36 => x_36_tb,
	x_37 => x_37_tb,
	x_38 => x_38_tb,
	x_39 => x_39_tb,
	x_40 => x_40_tb,
	x_41 => x_41_tb,
	x_42 => x_42_tb,
	x_43 => x_43_tb,
	x_44 => x_44_tb,
	x_45 => x_45_tb,
	x_46 => x_46_tb,
	x_47 => x_47_tb,
	x_48 => x_48_tb,
	x_49 => x_49_tb,
	x_50 => x_50_tb,
	x_51 => x_51_tb,
	x_52 => x_52_tb,
	x_53 => x_53_tb,
	x_54 => x_54_tb,
	x_55 => x_55_tb,
	x_56 => x_56_tb,
	x_57 => x_57_tb,
	x_58 => x_58_tb,
	x_59 => x_59_tb,
	x_60 => x_60_tb,
	x_61 => x_61_tb,
	x_62 => x_62_tb,
	x_63 => x_63_tb,
	x_64 => x_64_tb,
	x_65 => x_65_tb,
	x_66 => x_66_tb,
	x_67 => x_67_tb,
	x_68 => x_68_tb,
	x_69 => x_69_tb,
	x_70 => x_70_tb,
	x_71 => x_71_tb,
	x_72 => x_72_tb,
	x_73 => x_73_tb,
	x_74 => x_74_tb,
	x_75 => x_75_tb,
	x_76 => x_76_tb,
	x_77 => x_77_tb,
	x_78 => x_78_tb,
	x_79 => x_79_tb,
	x_80 => x_80_tb,
	x_81 => x_81_tb,
	x_82 => x_82_tb,
	x_83 => x_83_tb,
	x_84 => x_84_tb,
	x_85 => x_85_tb,
	x_86 => x_86_tb,
	x_87 => x_87_tb,
	x_88 => x_88_tb,
	x_89 => x_89_tb,
	x_90 => x_90_tb,
	x_91 => x_91_tb,
	x_92 => x_92_tb,
	x_93 => x_93_tb,
	x_94 => x_94_tb,
	x_95 => x_95_tb,
	x_96 => x_96_tb,
	x_97 => x_97_tb,
	x_98 => x_98_tb,
	x_99 => x_99_tb,
	x_100 => x_100_tb,
	x_101 => x_101_tb,
	x_102 => x_102_tb,
	x_103 => x_103_tb,
	x_104 => x_104_tb,
	x_105 => x_105_tb,
	x_106 => x_106_tb,
	x_107 => x_107_tb,
	x_108 => x_108_tb,
	x_109 => x_109_tb,
	x_110 => x_110_tb,
	x_111 => x_111_tb,
	x_112 => x_112_tb,
	x_113 => x_113_tb,
	x_114 => x_114_tb,
	x_115 => x_115_tb,
	x_116 => x_116_tb,
	x_117 => x_117_tb,
	x_118 => x_118_tb,
	x_119 => x_119_tb,
	x_120 => x_120_tb,
	x_121 => x_121_tb,
	x_122 => x_122_tb,
	x_123 => x_123_tb,
	x_124 => x_124_tb,
	x_125 => x_125_tb,
	x_126 => x_126_tb,
	x_127 => x_127_tb,
	x_128 => x_128_tb,
	x_129 => x_129_tb,
	x_130 => x_130_tb,
	x_131 => x_131_tb,
	x_132 => x_132_tb,
	x_133 => x_133_tb,
	x_134 => x_134_tb,
	x_135 => x_135_tb,
	x_136 => x_136_tb,
	x_137 => x_137_tb,
	x_138 => x_138_tb,
	x_139 => x_139_tb,
	x_140 => x_140_tb,
	x_141 => x_141_tb,
	x_142 => x_142_tb,
	x_143 => x_143_tb,
	x_144 => x_144_tb,
	x_145 => x_145_tb,
	x_146 => x_146_tb,
	x_147 => x_147_tb,
	x_148 => x_148_tb,
	x_149 => x_149_tb,
	x_150 => x_150_tb,
	x_151 => x_151_tb,
	x_152 => x_152_tb,
	x_153 => x_153_tb,
	x_154 => x_154_tb,
	x_155 => x_155_tb,
	x_156 => x_156_tb,
	x_157 => x_157_tb,
	x_158 => x_158_tb,
	x_159 => x_159_tb,
	x_160 => x_160_tb,
	x_161 => x_161_tb,
	x_162 => x_162_tb,
	x_163 => x_163_tb,
	x_164 => x_164_tb,
	x_165 => x_165_tb,
	x_166 => x_166_tb,
	x_167 => x_167_tb,
	x_168 => x_168_tb,
	x_169 => x_169_tb,
	x_170 => x_170_tb,
	x_171 => x_171_tb,
	x_172 => x_172_tb,
	x_173 => x_173_tb,
	x_174 => x_174_tb,
	x_175 => x_175_tb,
	x_176 => x_176_tb,
	x_177 => x_177_tb,
	x_178 => x_178_tb,
	x_179 => x_179_tb,
	x_180 => x_180_tb,
	x_181 => x_181_tb,
	x_182 => x_182_tb,
	x_183 => x_183_tb,
	x_184 => x_184_tb,
	x_185 => x_185_tb,
	x_186 => x_186_tb,
	x_187 => x_187_tb,
	x_188 => x_188_tb,
	x_189 => x_189_tb,
	x_190 => x_190_tb,
	x_191 => x_191_tb,
	x_192 => x_192_tb,
	x_193 => x_193_tb,
	x_194 => x_194_tb,
	x_195 => x_195_tb,
	x_196 => x_196_tb,
	x_197 => x_197_tb,
	x_198 => x_198_tb,
	x_199 => x_199_tb,
	x_200 => x_200_tb,
	x_201 => x_201_tb,
	x_202 => x_202_tb,
	x_203 => x_203_tb,
	x_204 => x_204_tb,
	x_205 => x_205_tb,
	x_206 => x_206_tb,
	x_207 => x_207_tb,
	x_208 => x_208_tb,
	x_209 => x_209_tb,
	x_210 => x_210_tb,
	x_211 => x_211_tb,
	x_212 => x_212_tb,
	x_213 => x_213_tb,
	x_214 => x_214_tb,
	x_215 => x_215_tb,
	x_216 => x_216_tb,
	x_217 => x_217_tb,
	x_218 => x_218_tb,
	x_219 => x_219_tb,
	x_220 => x_220_tb,
	x_221 => x_221_tb,
	x_222 => x_222_tb,
	x_223 => x_223_tb,
	x_224 => x_224_tb,
	x_225 => x_225_tb,
	x_226 => x_226_tb,
	x_227 => x_227_tb,
	x_228 => x_228_tb,
	x_229 => x_229_tb,
	x_230 => x_230_tb,
	x_231 => x_231_tb,
	x_232 => x_232_tb,
	x_233 => x_233_tb,
	x_234 => x_234_tb,
	x_235 => x_235_tb,
	x_236 => x_236_tb,
	x_237 => x_237_tb,
	x_238 => x_238_tb,
	x_239 => x_239_tb,
	x_240 => x_240_tb,
	x_241 => x_241_tb,
	x_242 => x_242_tb,
	x_243 => x_243_tb,
	x_244 => x_244_tb,
	x_245 => x_245_tb,
	x_246 => x_246_tb,
	x_247 => x_247_tb,
	x_248 => x_248_tb,
	x_249 => x_249_tb,
	x_250 => x_250_tb,
	x_251 => x_251_tb,
	x_252 => x_252_tb,
	x_253 => x_253_tb,
	x_254 => x_254_tb,
	x_255 => x_255_tb,
	x_256 => x_256_tb,
	x_257 => x_257_tb,
	x_258 => x_258_tb,
	x_259 => x_259_tb,
	x_260 => x_260_tb,
	x_261 => x_261_tb,
	x_262 => x_262_tb,
	x_263 => x_263_tb,
	x_264 => x_264_tb,
	x_265 => x_265_tb,
	x_266 => x_266_tb,
	x_267 => x_267_tb,
	x_268 => x_268_tb,
	x_269 => x_269_tb,
	x_270 => x_270_tb,
	x_271 => x_271_tb,
	x_272 => x_272_tb,
	x_273 => x_273_tb,
	x_274 => x_274_tb,
	x_275 => x_275_tb,
	x_276 => x_276_tb,
	x_277 => x_277_tb,
	x_278 => x_278_tb,
	x_279 => x_279_tb,
	x_280 => x_280_tb,
	x_281 => x_281_tb,
	x_282 => x_282_tb,
	x_283 => x_283_tb,
	x_284 => x_284_tb,
	x_285 => x_285_tb,
	x_286 => x_286_tb,
	x_287 => x_287_tb,
	x_288 => x_288_tb,
	x_289 => x_289_tb,
	x_290 => x_290_tb,
	x_291 => x_291_tb,
	x_292 => x_292_tb,
	x_293 => x_293_tb,
	x_294 => x_294_tb,
	x_295 => x_295_tb,
	x_296 => x_296_tb,
	x_297 => x_297_tb,
	x_298 => x_298_tb,
	x_299 => x_299_tb,
	x_300 => x_300_tb,
	x_301 => x_301_tb,
	x_302 => x_302_tb,
	x_303 => x_303_tb,
	x_304 => x_304_tb,
	x_305 => x_305_tb,
	x_306 => x_306_tb,
	x_307 => x_307_tb,
	x_308 => x_308_tb,
	x_309 => x_309_tb,
	x_310 => x_310_tb,
	x_311 => x_311_tb,
	x_312 => x_312_tb,
	x_313 => x_313_tb,
	x_314 => x_314_tb,
	x_315 => x_315_tb,
	x_316 => x_316_tb,
	x_317 => x_317_tb,
	x_318 => x_318_tb,
	x_319 => x_319_tb,
	x_320 => x_320_tb,
	x_321 => x_321_tb,
	x_322 => x_322_tb,
	x_323 => x_323_tb,
	x_324 => x_324_tb,
	x_325 => x_325_tb,
	x_326 => x_326_tb,
	x_327 => x_327_tb,
	x_328 => x_328_tb,
	x_329 => x_329_tb,
	x_330 => x_330_tb,
	x_331 => x_331_tb,
	x_332 => x_332_tb,
	x_333 => x_333_tb,
	x_334 => x_334_tb,
	x_335 => x_335_tb,
	x_336 => x_336_tb,
	x_337 => x_337_tb,
	x_338 => x_338_tb,
	x_339 => x_339_tb,
	x_340 => x_340_tb,
	x_341 => x_341_tb,
	x_342 => x_342_tb,
	x_343 => x_343_tb,
	x_344 => x_344_tb,
	x_345 => x_345_tb,
	x_346 => x_346_tb,
	x_347 => x_347_tb,
	x_348 => x_348_tb,
	x_349 => x_349_tb,
	x_350 => x_350_tb,
	x_351 => x_351_tb,
	x_352 => x_352_tb,
	x_353 => x_353_tb,
	x_354 => x_354_tb,
	x_355 => x_355_tb,
	x_356 => x_356_tb,
	x_357 => x_357_tb,
	x_358 => x_358_tb,
	x_359 => x_359_tb,
	x_360 => x_360_tb,
	x_361 => x_361_tb,
	x_362 => x_362_tb,
	x_363 => x_363_tb,
	x_364 => x_364_tb,
	x_365 => x_365_tb,
	x_366 => x_366_tb,
	x_367 => x_367_tb,
	x_368 => x_368_tb,
	x_369 => x_369_tb,
	x_370 => x_370_tb,
	x_371 => x_371_tb,
	x_372 => x_372_tb,
	x_373 => x_373_tb,
	x_374 => x_374_tb,
	x_375 => x_375_tb,
	x_376 => x_376_tb,
	x_377 => x_377_tb,
	x_378 => x_378_tb,
	x_379 => x_379_tb,
	x_380 => x_380_tb,
	x_381 => x_381_tb,
	x_382 => x_382_tb,
	x_383 => x_383_tb,
	x_384 => x_384_tb,
	x_385 => x_385_tb,
	x_386 => x_386_tb,
	x_387 => x_387_tb,
	x_388 => x_388_tb,
	x_389 => x_389_tb,
	x_390 => x_390_tb,
	x_391 => x_391_tb,
	x_392 => x_392_tb,
	x_393 => x_393_tb,
	x_394 => x_394_tb,
	x_395 => x_395_tb,
	x_396 => x_396_tb,
	x_397 => x_397_tb,
	x_398 => x_398_tb,
	x_399 => x_399_tb,
	x_400 => x_400_tb,
	x_401 => x_401_tb,
	x_402 => x_402_tb,
	x_403 => x_403_tb,
	x_404 => x_404_tb,
	x_405 => x_405_tb,
	x_406 => x_406_tb,
	x_407 => x_407_tb,
	x_408 => x_408_tb,
	x_409 => x_409_tb,
	x_410 => x_410_tb,
	x_411 => x_411_tb,
	x_412 => x_412_tb,
	x_413 => x_413_tb,
	x_414 => x_414_tb,
	x_415 => x_415_tb,
	x_416 => x_416_tb,
	x_417 => x_417_tb,
	x_418 => x_418_tb,
	x_419 => x_419_tb,
	x_420 => x_420_tb,
	x_421 => x_421_tb,
	x_422 => x_422_tb,
	x_423 => x_423_tb,
	x_424 => x_424_tb,
	x_425 => x_425_tb,
	x_426 => x_426_tb,
	x_427 => x_427_tb,
	x_428 => x_428_tb,
	x_429 => x_429_tb,
	x_430 => x_430_tb,
	x_431 => x_431_tb,
	x_432 => x_432_tb,
	x_433 => x_433_tb,
	x_434 => x_434_tb,
	x_435 => x_435_tb,
	x_436 => x_436_tb,
	x_437 => x_437_tb,
	x_438 => x_438_tb,
	x_439 => x_439_tb,
	x_440 => x_440_tb,
	x_441 => x_441_tb,
	x_442 => x_442_tb,
	x_443 => x_443_tb,
	x_444 => x_444_tb,
	x_445 => x_445_tb,
	x_446 => x_446_tb,
	x_447 => x_447_tb,
	x_448 => x_448_tb,
	x_449 => x_449_tb,
	x_450 => x_450_tb,
	x_451 => x_451_tb,
	x_452 => x_452_tb,
	x_453 => x_453_tb,
	x_454 => x_454_tb,
	x_455 => x_455_tb,
	x_456 => x_456_tb,
	x_457 => x_457_tb,
	x_458 => x_458_tb,
	x_459 => x_459_tb,
	x_460 => x_460_tb,
	x_461 => x_461_tb,
	x_462 => x_462_tb,
	x_463 => x_463_tb,
	x_464 => x_464_tb,
	x_465 => x_465_tb,
	x_466 => x_466_tb,
	x_467 => x_467_tb,
	x_468 => x_468_tb,
	x_469 => x_469_tb,
	x_470 => x_470_tb,
	x_471 => x_471_tb,
	x_472 => x_472_tb,
	x_473 => x_473_tb,
	x_474 => x_474_tb,
	x_475 => x_475_tb,
	x_476 => x_476_tb,
	x_477 => x_477_tb,
	x_478 => x_478_tb,
	x_479 => x_479_tb,
	x_480 => x_480_tb,
	x_481 => x_481_tb,
	x_482 => x_482_tb,
	x_483 => x_483_tb,
	x_484 => x_484_tb,
	x_485 => x_485_tb,
	x_486 => x_486_tb,
	x_487 => x_487_tb,
	x_488 => x_488_tb,
	x_489 => x_489_tb,
	x_490 => x_490_tb,
	x_491 => x_491_tb,
	x_492 => x_492_tb,
	x_493 => x_493_tb,
	x_494 => x_494_tb,
	x_495 => x_495_tb,
	x_496 => x_496_tb,
	x_497 => x_497_tb,
	x_498 => x_498_tb,
	x_499 => x_499_tb,
	x_500 => x_500_tb,
	x_501 => x_501_tb,
	x_502 => x_502_tb,
	x_503 => x_503_tb,
	x_504 => x_504_tb,
	x_505 => x_505_tb,
	x_506 => x_506_tb,
	x_507 => x_507_tb,
	x_508 => x_508_tb,
	x_509 => x_509_tb,
	x_510 => x_510_tb,
	x_511 => x_511_tb,
	x_512 => x_512_tb,
	x_513 => x_513_tb,
	x_514 => x_514_tb,
	x_515 => x_515_tb,
	x_516 => x_516_tb,
	x_517 => x_517_tb,
	x_518 => x_518_tb,
	x_519 => x_519_tb,
	x_520 => x_520_tb,
	x_521 => x_521_tb,
	x_522 => x_522_tb,
	x_523 => x_523_tb,
	x_524 => x_524_tb,
	x_525 => x_525_tb,
	x_526 => x_526_tb,
	x_527 => x_527_tb,
	x_528 => x_528_tb,
	x_529 => x_529_tb,
	x_530 => x_530_tb,
	x_531 => x_531_tb,
	x_532 => x_532_tb,
	x_533 => x_533_tb,
	x_534 => x_534_tb,
	x_535 => x_535_tb,
	x_536 => x_536_tb,
	x_537 => x_537_tb,
	x_538 => x_538_tb,
	x_539 => x_539_tb,
	x_540 => x_540_tb,
	x_541 => x_541_tb,
	x_542 => x_542_tb,
	x_543 => x_543_tb,
	x_544 => x_544_tb,
	x_545 => x_545_tb,
	x_546 => x_546_tb,
	x_547 => x_547_tb,
	x_548 => x_548_tb,
	x_549 => x_549_tb,
	x_550 => x_550_tb,
	x_551 => x_551_tb,
	x_552 => x_552_tb,
	x_553 => x_553_tb,
	x_554 => x_554_tb,
	x_555 => x_555_tb,
	x_556 => x_556_tb,
	x_557 => x_557_tb,
	x_558 => x_558_tb,
	x_559 => x_559_tb,
	x_560 => x_560_tb,
	x_561 => x_561_tb,
	x_562 => x_562_tb,
	x_563 => x_563_tb,
	x_564 => x_564_tb,
	x_565 => x_565_tb,
	x_566 => x_566_tb,
	x_567 => x_567_tb,
	x_568 => x_568_tb,
	x_569 => x_569_tb,
	x_570 => x_570_tb,
	x_571 => x_571_tb,
	x_572 => x_572_tb,
	x_573 => x_573_tb,
	x_574 => x_574_tb,
	x_575 => x_575_tb,
	x_576 => x_576_tb,
	x_577 => x_577_tb,
	x_578 => x_578_tb,
	x_579 => x_579_tb,
	x_580 => x_580_tb,
	x_581 => x_581_tb,
	x_582 => x_582_tb,
	x_583 => x_583_tb,
	x_584 => x_584_tb,
	x_585 => x_585_tb,
	x_586 => x_586_tb,
	x_587 => x_587_tb,
	x_588 => x_588_tb,
	x_589 => x_589_tb,
	x_590 => x_590_tb,
	x_591 => x_591_tb,
	x_592 => x_592_tb,
	x_593 => x_593_tb,
	x_594 => x_594_tb,
	x_595 => x_595_tb,
	x_596 => x_596_tb,
	x_597 => x_597_tb,
	x_598 => x_598_tb,
	x_599 => x_599_tb,
	x_600 => x_600_tb,
	x_601 => x_601_tb,
	x_602 => x_602_tb,
	x_603 => x_603_tb,
	x_604 => x_604_tb,
	x_605 => x_605_tb,
	x_606 => x_606_tb,
	x_607 => x_607_tb,
	x_608 => x_608_tb,
	x_609 => x_609_tb,
	x_610 => x_610_tb,
	x_611 => x_611_tb,
	x_612 => x_612_tb,
	x_613 => x_613_tb,
	x_614 => x_614_tb,
	x_615 => x_615_tb,
	x_616 => x_616_tb,
	x_617 => x_617_tb,
	x_618 => x_618_tb,
	x_619 => x_619_tb,
	x_620 => x_620_tb,
	x_621 => x_621_tb,
	x_622 => x_622_tb,
	x_623 => x_623_tb,
	x_624 => x_624_tb,
	x_625 => x_625_tb,
	x_626 => x_626_tb,
	x_627 => x_627_tb,
	x_628 => x_628_tb,
	x_629 => x_629_tb,
	x_630 => x_630_tb,
	x_631 => x_631_tb,
	x_632 => x_632_tb,
	x_633 => x_633_tb,
	x_634 => x_634_tb,
	x_635 => x_635_tb,
	x_636 => x_636_tb,
	x_637 => x_637_tb,
	x_638 => x_638_tb,
	x_639 => x_639_tb,
	x_640 => x_640_tb,
	x_641 => x_641_tb,
	x_642 => x_642_tb,
	x_643 => x_643_tb,
	x_644 => x_644_tb,
	x_645 => x_645_tb,
	x_646 => x_646_tb,
	x_647 => x_647_tb,
	x_648 => x_648_tb,
	x_649 => x_649_tb,
	x_650 => x_650_tb,
	x_651 => x_651_tb,
	x_652 => x_652_tb,
	x_653 => x_653_tb,
	x_654 => x_654_tb,
	x_655 => x_655_tb,
	x_656 => x_656_tb,
	x_657 => x_657_tb,
	x_658 => x_658_tb,
	x_659 => x_659_tb,
	x_660 => x_660_tb,
	x_661 => x_661_tb,
	x_662 => x_662_tb,
	x_663 => x_663_tb,
	x_664 => x_664_tb,
	x_665 => x_665_tb,
	x_666 => x_666_tb,
	x_667 => x_667_tb,
	x_668 => x_668_tb,
	x_669 => x_669_tb,
	x_670 => x_670_tb,
	x_671 => x_671_tb,
	x_672 => x_672_tb,
	x_673 => x_673_tb,
	x_674 => x_674_tb,
	x_675 => x_675_tb,
	x_676 => x_676_tb,
	x_677 => x_677_tb,
	x_678 => x_678_tb,
	x_679 => x_679_tb,
	x_680 => x_680_tb,
	x_681 => x_681_tb,
	x_682 => x_682_tb,
	x_683 => x_683_tb,
	x_684 => x_684_tb,
	x_685 => x_685_tb,
	x_686 => x_686_tb,
	x_687 => x_687_tb,
	x_688 => x_688_tb,
	x_689 => x_689_tb,
	x_690 => x_690_tb,
	x_691 => x_691_tb,
	x_692 => x_692_tb,
	x_693 => x_693_tb,
	x_694 => x_694_tb,
	x_695 => x_695_tb,
	x_696 => x_696_tb,
	x_697 => x_697_tb,
	x_698 => x_698_tb,
	x_699 => x_699_tb,
	x_700 => x_700_tb,
	x_701 => x_701_tb,
	x_702 => x_702_tb,
	x_703 => x_703_tb,
	x_704 => x_704_tb,
	x_705 => x_705_tb,
	x_706 => x_706_tb,
	x_707 => x_707_tb,
	x_708 => x_708_tb,
	x_709 => x_709_tb,
	x_710 => x_710_tb,
	x_711 => x_711_tb,
	x_712 => x_712_tb,
	x_713 => x_713_tb,
	x_714 => x_714_tb,
	x_715 => x_715_tb,
	x_716 => x_716_tb,
	x_717 => x_717_tb,
	x_718 => x_718_tb,
	x_719 => x_719_tb,
	x_720 => x_720_tb,
	x_721 => x_721_tb,
	x_722 => x_722_tb,
	x_723 => x_723_tb,
	x_724 => x_724_tb,
	x_725 => x_725_tb,
	x_726 => x_726_tb,
	x_727 => x_727_tb,
	x_728 => x_728_tb,
	x_729 => x_729_tb,
	x_730 => x_730_tb,
	x_731 => x_731_tb,
	x_732 => x_732_tb,
	x_733 => x_733_tb,
	x_734 => x_734_tb,
	x_735 => x_735_tb,
	x_736 => x_736_tb,
	x_737 => x_737_tb,
	x_738 => x_738_tb,
	x_739 => x_739_tb,
	x_740 => x_740_tb,
	x_741 => x_741_tb,
	x_742 => x_742_tb,
	x_743 => x_743_tb,
	x_744 => x_744_tb,
	x_745 => x_745_tb,
	x_746 => x_746_tb,
	x_747 => x_747_tb,
	x_748 => x_748_tb,
	x_749 => x_749_tb,
	x_750 => x_750_tb,
	x_751 => x_751_tb,
	x_752 => x_752_tb,
	x_753 => x_753_tb,
	x_754 => x_754_tb,
	x_755 => x_755_tb,
	x_756 => x_756_tb,
	x_757 => x_757_tb,
	x_758 => x_758_tb,
	x_759 => x_759_tb,
	x_760 => x_760_tb,
	x_761 => x_761_tb,
	x_762 => x_762_tb,
	x_763 => x_763_tb,
	x_764 => x_764_tb,
	x_765 => x_765_tb,
	x_766 => x_766_tb,
	x_767 => x_767_tb,
	x_768 => x_768_tb,
	x_769 => x_769_tb,
	x_770 => x_770_tb,
	x_771 => x_771_tb,
	x_772 => x_772_tb,
	x_773 => x_773_tb,
	x_774 => x_774_tb,
	x_775 => x_775_tb,
	x_776 => x_776_tb,
	x_777 => x_777_tb,
	x_778 => x_778_tb,
	x_779 => x_779_tb,
	x_780 => x_780_tb,
	x_781 => x_781_tb,
	x_782 => x_782_tb,
	x_783 => x_783_tb,
	y => y_tb
    );
clk_process: process
   begin
       while now < 1000 ns loop
       clk_tb <= '0';
       wait for CLK_PERIOD / 2;
       clk_tb <= '1';
       wait for CLK_PERIOD / 2;
   end loop;
   wait;
end process;
stim_proc: process
   begin
       x_0_tb <= "0000000000000000"; 
       x_1_tb <= "0000000000000000"; 
       x_2_tb <= "0000000000000000"; 
       x_3_tb <= "0000000000000000"; 
       x_4_tb <= "0000000000000000"; 
       x_5_tb <= "0000000000000000"; 
       x_6_tb <= "0000000000000000"; 
       x_7_tb <= "0000000000000000"; 
       x_8_tb <= "0000000000000000"; 
       x_9_tb <= "0000000000000000"; 
       x_10_tb <= "0000000000000000"; 
       x_11_tb <= "0000000000000000"; 
       x_12_tb <= "0000000000000000"; 
       x_13_tb <= "0000000000000000"; 
       x_14_tb <= "0000000000000000"; 
       x_15_tb <= "0000000000000000"; 
       x_16_tb <= "0000000000000000"; 
       x_17_tb <= "0000000000000000"; 
       x_18_tb <= "0000000000000000"; 
       x_19_tb <= "0000000000000000"; 
       x_20_tb <= "0000000000000000"; 
       x_21_tb <= "0000000000000000"; 
       x_22_tb <= "0000000000000000"; 
       x_23_tb <= "0000000000000000"; 
       x_24_tb <= "0000000000000000"; 
       x_25_tb <= "0000000000000000"; 
       x_26_tb <= "0000000000000000"; 
       x_27_tb <= "0000000000000000"; 
       x_28_tb <= "0000000000000000"; 
       x_29_tb <= "0000000000000000"; 
       x_30_tb <= "0000000000000000"; 
       x_31_tb <= "0000000000000000"; 
       x_32_tb <= "0000000000000000"; 
       x_33_tb <= "0000000000000000"; 
       x_34_tb <= "0000000000000000"; 
       x_35_tb <= "0000000000000000"; 
       x_36_tb <= "0000000000000000"; 
       x_37_tb <= "0000000000000000"; 
       x_38_tb <= "0000000000000000"; 
       x_39_tb <= "0000000000000000"; 
       x_40_tb <= "0000000000000000"; 
       x_41_tb <= "0000000000000000"; 
       x_42_tb <= "0000000000000000"; 
       x_43_tb <= "0000000000000000"; 
       x_44_tb <= "0000000000000000"; 
       x_45_tb <= "0000000000000000"; 
       x_46_tb <= "0000000000000000"; 
       x_47_tb <= "0000000000000000"; 
       x_48_tb <= "0000000000000000"; 
       x_49_tb <= "0000000000000000"; 
       x_50_tb <= "0000000000000000"; 
       x_51_tb <= "0000000000000000"; 
       x_52_tb <= "0000000000000000"; 
       x_53_tb <= "0000000000000000"; 
       x_54_tb <= "0000000000000000"; 
       x_55_tb <= "0000000000000000"; 
       x_56_tb <= "0000000000000000"; 
       x_57_tb <= "0000000000000000"; 
       x_58_tb <= "0000000000000000"; 
       x_59_tb <= "0000000000000000"; 
       x_60_tb <= "0000000000000000"; 
       x_61_tb <= "0000000000000000"; 
       x_62_tb <= "0000000000000000"; 
       x_63_tb <= "0000000000000000"; 
       x_64_tb <= "0000000000000000"; 
       x_65_tb <= "0000000000000000"; 
       x_66_tb <= "0000000000000000"; 
       x_67_tb <= "0000000000000000"; 
       x_68_tb <= "0000000000000000"; 
       x_69_tb <= "0000000000000000"; 
       x_70_tb <= "0000000000000000"; 
       x_71_tb <= "0000000000000000"; 
       x_72_tb <= "0000000000000000"; 
       x_73_tb <= "0000000000000000"; 
       x_74_tb <= "0000000000000000"; 
       x_75_tb <= "0000000000000000"; 
       x_76_tb <= "0000000000000000"; 
       x_77_tb <= "0000000000000000"; 
       x_78_tb <= "0000000000000000"; 
       x_79_tb <= "0000000000000000"; 
       x_80_tb <= "0000000000000000"; 
       x_81_tb <= "0000000000000000"; 
       x_82_tb <= "0000000000000000"; 
       x_83_tb <= "0000000000000000"; 
       x_84_tb <= "0000000000000000"; 
       x_85_tb <= "0000000000000000"; 
       x_86_tb <= "0000000000000000"; 
       x_87_tb <= "0000000000000000"; 
       x_88_tb <= "0000000000000000"; 
       x_89_tb <= "0000000000000000"; 
       x_90_tb <= "0000000000000000"; 
       x_91_tb <= "0000000000000000"; 
       x_92_tb <= "0000000000000000"; 
       x_93_tb <= "0000000000000000"; 
       x_94_tb <= "0000000000000000"; 
       x_95_tb <= "0000000000000000"; 
       x_96_tb <= "0000000000000000"; 
       x_97_tb <= "0000000000000000"; 
       x_98_tb <= "0000000000000000"; 
       x_99_tb <= "0000000000000000"; 
       x_100_tb <= "0000000000000000"; 
       x_101_tb <= "0000000000000000"; 
       x_102_tb <= "0000000000000000"; 
       x_103_tb <= "0000000000000000"; 
       x_104_tb <= "0000000000000000"; 
       x_105_tb <= "0000000000000000"; 
       x_106_tb <= "0000000000000000"; 
       x_107_tb <= "0000000000000000"; 
       x_108_tb <= "0000000000000000"; 
       x_109_tb <= "0000000000000000"; 
       x_110_tb <= "0000000000000000"; 
       x_111_tb <= "0000000000000000"; 
       x_112_tb <= "0000000000000000"; 
       x_113_tb <= "0000000000000000"; 
       x_114_tb <= "0000000000000000"; 
       x_115_tb <= "0000000000000000"; 
       x_116_tb <= "0000000000000000"; 
       x_117_tb <= "0000000000000000"; 
       x_118_tb <= "0000000000000000"; 
       x_119_tb <= "0000000000000000"; 
       x_120_tb <= "0000000000000000"; 
       x_121_tb <= "0000000000000000"; 
       x_122_tb <= "0000000000000000"; 
       x_123_tb <= "0000000000000000"; 
       x_124_tb <= "0000000011001000"; 
       x_125_tb <= "0000000011111110"; 
       x_126_tb <= "0000000000000000"; 
       x_127_tb <= "0000000000000000"; 
       x_128_tb <= "0000000000000000"; 
       x_129_tb <= "0000000000000000"; 
       x_130_tb <= "0000000000000000"; 
       x_131_tb <= "0000000000000000"; 
       x_132_tb <= "0000000000000000"; 
       x_133_tb <= "0000000000000000"; 
       x_134_tb <= "0000000000000000"; 
       x_135_tb <= "0000000000000000"; 
       x_136_tb <= "0000000000000000"; 
       x_137_tb <= "0000000000000000"; 
       x_138_tb <= "0000000000000000"; 
       x_139_tb <= "0000000000000000"; 
       x_140_tb <= "0000000000000000"; 
       x_141_tb <= "0000000000000000"; 
       x_142_tb <= "0000000000000000"; 
       x_143_tb <= "0000000000000000"; 
       x_144_tb <= "0000000000000000"; 
       x_145_tb <= "0000000000000000"; 
       x_146_tb <= "0000000000000000"; 
       x_147_tb <= "0000000000000000"; 
       x_148_tb <= "0000000000000000"; 
       x_149_tb <= "0000000000000000"; 
       x_150_tb <= "0000000000000000"; 
       x_151_tb <= "0000000000000000"; 
       x_152_tb <= "0000000011010100"; 
       x_153_tb <= "0000000011111101"; 
       x_154_tb <= "0000000000000000"; 
       x_155_tb <= "0000000000000000"; 
       x_156_tb <= "0000000000000000"; 
       x_157_tb <= "0000000000000000"; 
       x_158_tb <= "0000000000000000"; 
       x_159_tb <= "0000000000000000"; 
       x_160_tb <= "0000000000000000"; 
       x_161_tb <= "0000000000000000"; 
       x_162_tb <= "0000000000000000"; 
       x_163_tb <= "0000000000000000"; 
       x_164_tb <= "0000000000000000"; 
       x_165_tb <= "0000000000000000"; 
       x_166_tb <= "0000000000000000"; 
       x_167_tb <= "0000000000000000"; 
       x_168_tb <= "0000000000000000"; 
       x_169_tb <= "0000000000000000"; 
       x_170_tb <= "0000000000000000"; 
       x_171_tb <= "0000000000000000"; 
       x_172_tb <= "0000000000000000"; 
       x_173_tb <= "0000000000000000"; 
       x_174_tb <= "0000000000000000"; 
       x_175_tb <= "0000000000000000"; 
       x_176_tb <= "0000000000000000"; 
       x_177_tb <= "0000000000000000"; 
       x_178_tb <= "0000000000000000"; 
       x_179_tb <= "0000000000000000"; 
       x_180_tb <= "0000000010100110"; 
       x_181_tb <= "0000000011111101"; 
       x_182_tb <= "0000000000000000"; 
       x_183_tb <= "0000000000000000"; 
       x_184_tb <= "0000000000000000"; 
       x_185_tb <= "0000000000000000"; 
       x_186_tb <= "0000000000000000"; 
       x_187_tb <= "0000000000000000"; 
       x_188_tb <= "0000000000000000"; 
       x_189_tb <= "0000000000000000"; 
       x_190_tb <= "0000000000000000"; 
       x_191_tb <= "0000000000000000"; 
       x_192_tb <= "0000000000000000"; 
       x_193_tb <= "0000000000000000"; 
       x_194_tb <= "0000000000000000"; 
       x_195_tb <= "0000000000000000"; 
       x_196_tb <= "0000000000000000"; 
       x_197_tb <= "0000000000000000"; 
       x_198_tb <= "0000000000000000"; 
       x_199_tb <= "0000000000000000"; 
       x_200_tb <= "0000000000000000"; 
       x_201_tb <= "0000000000000000"; 
       x_202_tb <= "0000000000000000"; 
       x_203_tb <= "0000000000000000"; 
       x_204_tb <= "0000000000000000"; 
       x_205_tb <= "0000000000000000"; 
       x_206_tb <= "0000000000000000"; 
       x_207_tb <= "0000000010010010"; 
       x_208_tb <= "0000000011111011"; 
       x_209_tb <= "0000000011111101"; 
       x_210_tb <= "0000000010000000"; 
       x_211_tb <= "0000000000000000"; 
       x_212_tb <= "0000000000000000"; 
       x_213_tb <= "0000000000000000"; 
       x_214_tb <= "0000000000000000"; 
       x_215_tb <= "0000000000000000"; 
       x_216_tb <= "0000000000000000"; 
       x_217_tb <= "0000000000000000"; 
       x_218_tb <= "0000000000000000"; 
       x_219_tb <= "0000000000000000"; 
       x_220_tb <= "0000000000000000"; 
       x_221_tb <= "0000000000000000"; 
       x_222_tb <= "0000000000000000"; 
       x_223_tb <= "0000000000000000"; 
       x_224_tb <= "0000000000000000"; 
       x_225_tb <= "0000000000000000"; 
       x_226_tb <= "0000000000000000"; 
       x_227_tb <= "0000000000000000"; 
       x_228_tb <= "0000000000000000"; 
       x_229_tb <= "0000000000000000"; 
       x_230_tb <= "0000000000000000"; 
       x_231_tb <= "0000000000000000"; 
       x_232_tb <= "0000000000000000"; 
       x_233_tb <= "0000000000000000"; 
       x_234_tb <= "0000000000000000"; 
       x_235_tb <= "0000000011000000"; 
       x_236_tb <= "0000000011110101"; 
       x_237_tb <= "0000000011111101"; 
       x_238_tb <= "0000000011000100"; 
       x_239_tb <= "0000000000000000"; 
       x_240_tb <= "0000000000000000"; 
       x_241_tb <= "0000000000000000"; 
       x_242_tb <= "0000000000000000"; 
       x_243_tb <= "0000000000000000"; 
       x_244_tb <= "0000000000000000"; 
       x_245_tb <= "0000000000000000"; 
       x_246_tb <= "0000000000000000"; 
       x_247_tb <= "0000000000000000"; 
       x_248_tb <= "0000000000000000"; 
       x_249_tb <= "0000000000000000"; 
       x_250_tb <= "0000000000000000"; 
       x_251_tb <= "0000000000000000"; 
       x_252_tb <= "0000000000000000"; 
       x_253_tb <= "0000000000000000"; 
       x_254_tb <= "0000000000000000"; 
       x_255_tb <= "0000000000000000"; 
       x_256_tb <= "0000000000000000"; 
       x_257_tb <= "0000000000000000"; 
       x_258_tb <= "0000000000000000"; 
       x_259_tb <= "0000000000000000"; 
       x_260_tb <= "0000000000000000"; 
       x_261_tb <= "0000000000000000"; 
       x_262_tb <= "0000000000000000"; 
       x_263_tb <= "0000000000000000"; 
       x_264_tb <= "0000000011101011"; 
       x_265_tb <= "0000000011111110"; 
       x_266_tb <= "0000000011000100"; 
       x_267_tb <= "0000000000000000"; 
       x_268_tb <= "0000000000000000"; 
       x_269_tb <= "0000000000000000"; 
       x_270_tb <= "0000000000000000"; 
       x_271_tb <= "0000000000000000"; 
       x_272_tb <= "0000000000000000"; 
       x_273_tb <= "0000000000000000"; 
       x_274_tb <= "0000000000000000"; 
       x_275_tb <= "0000000000000000"; 
       x_276_tb <= "0000000000000000"; 
       x_277_tb <= "0000000000000000"; 
       x_278_tb <= "0000000000000000"; 
       x_279_tb <= "0000000000000000"; 
       x_280_tb <= "0000000000000000"; 
       x_281_tb <= "0000000000000000"; 
       x_282_tb <= "0000000000000000"; 
       x_283_tb <= "0000000000000000"; 
       x_284_tb <= "0000000000000000"; 
       x_285_tb <= "0000000000000000"; 
       x_286_tb <= "0000000000000000"; 
       x_287_tb <= "0000000000000000"; 
       x_288_tb <= "0000000000000000"; 
       x_289_tb <= "0000000000000000"; 
       x_290_tb <= "0000000000000000"; 
       x_291_tb <= "0000000000000000"; 
       x_292_tb <= "0000000010010111"; 
       x_293_tb <= "0000000011111101"; 
       x_294_tb <= "0000000011011110"; 
       x_295_tb <= "0000000010010000"; 
       x_296_tb <= "0000000000000000"; 
       x_297_tb <= "0000000000000000"; 
       x_298_tb <= "0000000000000000"; 
       x_299_tb <= "0000000000000000"; 
       x_300_tb <= "0000000000000000"; 
       x_301_tb <= "0000000000000000"; 
       x_302_tb <= "0000000000000000"; 
       x_303_tb <= "0000000000000000"; 
       x_304_tb <= "0000000000000000"; 
       x_305_tb <= "0000000000000000"; 
       x_306_tb <= "0000000000000000"; 
       x_307_tb <= "0000000000000000"; 
       x_308_tb <= "0000000000000000"; 
       x_309_tb <= "0000000000000000"; 
       x_310_tb <= "0000000000000000"; 
       x_311_tb <= "0000000000000000"; 
       x_312_tb <= "0000000000000000"; 
       x_313_tb <= "0000000000000000"; 
       x_314_tb <= "0000000000000000"; 
       x_315_tb <= "0000000000000000"; 
       x_316_tb <= "0000000000000000"; 
       x_317_tb <= "0000000000000000"; 
       x_318_tb <= "0000000000000000"; 
       x_319_tb <= "0000000000000000"; 
       x_320_tb <= "0000000010001010"; 
       x_321_tb <= "0000000011111101"; 
       x_322_tb <= "0000000011101011"; 
       x_323_tb <= "0000000011011000"; 
       x_324_tb <= "0000000000000000"; 
       x_325_tb <= "0000000000000000"; 
       x_326_tb <= "0000000000000000"; 
       x_327_tb <= "0000000000000000"; 
       x_328_tb <= "0000000000000000"; 
       x_329_tb <= "0000000000000000"; 
       x_330_tb <= "0000000000000000"; 
       x_331_tb <= "0000000000000000"; 
       x_332_tb <= "0000000000000000"; 
       x_333_tb <= "0000000000000000"; 
       x_334_tb <= "0000000000000000"; 
       x_335_tb <= "0000000000000000"; 
       x_336_tb <= "0000000000000000"; 
       x_337_tb <= "0000000000000000"; 
       x_338_tb <= "0000000000000000"; 
       x_339_tb <= "0000000000000000"; 
       x_340_tb <= "0000000000000000"; 
       x_341_tb <= "0000000000000000"; 
       x_342_tb <= "0000000000000000"; 
       x_343_tb <= "0000000000000000"; 
       x_344_tb <= "0000000000000000"; 
       x_345_tb <= "0000000000000000"; 
       x_346_tb <= "0000000000000000"; 
       x_347_tb <= "0000000000000000"; 
       x_348_tb <= "0000000010100000"; 
       x_349_tb <= "0000000011111101"; 
       x_350_tb <= "0000000011100011"; 
       x_351_tb <= "0000000010101000"; 
       x_352_tb <= "0000000000000000"; 
       x_353_tb <= "0000000000000000"; 
       x_354_tb <= "0000000000000000"; 
       x_355_tb <= "0000000000000000"; 
       x_356_tb <= "0000000000000000"; 
       x_357_tb <= "0000000000000000"; 
       x_358_tb <= "0000000000000000"; 
       x_359_tb <= "0000000000000000"; 
       x_360_tb <= "0000000000000000"; 
       x_361_tb <= "0000000000000000"; 
       x_362_tb <= "0000000000000000"; 
       x_363_tb <= "0000000000000000"; 
       x_364_tb <= "0000000000000000"; 
       x_365_tb <= "0000000000000000"; 
       x_366_tb <= "0000000000000000"; 
       x_367_tb <= "0000000000000000"; 
       x_368_tb <= "0000000000000000"; 
       x_369_tb <= "0000000000000000"; 
       x_370_tb <= "0000000000000000"; 
       x_371_tb <= "0000000000000000"; 
       x_372_tb <= "0000000000000000"; 
       x_373_tb <= "0000000000000000"; 
       x_374_tb <= "0000000000000000"; 
       x_375_tb <= "0000000000000000"; 
       x_376_tb <= "0000000010100000"; 
       x_377_tb <= "0000000011111101"; 
       x_378_tb <= "0000000011111110"; 
       x_379_tb <= "0000000010011100"; 
       x_380_tb <= "0000000000000000"; 
       x_381_tb <= "0000000000000000"; 
       x_382_tb <= "0000000000000000"; 
       x_383_tb <= "0000000000000000"; 
       x_384_tb <= "0000000000000000"; 
       x_385_tb <= "0000000000000000"; 
       x_386_tb <= "0000000000000000"; 
       x_387_tb <= "0000000000000000"; 
       x_388_tb <= "0000000000000000"; 
       x_389_tb <= "0000000000000000"; 
       x_390_tb <= "0000000000000000"; 
       x_391_tb <= "0000000000000000"; 
       x_392_tb <= "0000000000000000"; 
       x_393_tb <= "0000000000000000"; 
       x_394_tb <= "0000000000000000"; 
       x_395_tb <= "0000000000000000"; 
       x_396_tb <= "0000000000000000"; 
       x_397_tb <= "0000000000000000"; 
       x_398_tb <= "0000000000000000"; 
       x_399_tb <= "0000000000000000"; 
       x_400_tb <= "0000000000000000"; 
       x_401_tb <= "0000000000000000"; 
       x_402_tb <= "0000000000000000"; 
       x_403_tb <= "0000000000000000"; 
       x_404_tb <= "0000000011111000"; 
       x_405_tb <= "0000000011110000"; 
       x_406_tb <= "0000000011111111"; 
       x_407_tb <= "0000000010011100"; 
       x_408_tb <= "0000000000000000"; 
       x_409_tb <= "0000000000000000"; 
       x_410_tb <= "0000000000000000"; 
       x_411_tb <= "0000000000000000"; 
       x_412_tb <= "0000000000000000"; 
       x_413_tb <= "0000000000000000"; 
       x_414_tb <= "0000000000000000"; 
       x_415_tb <= "0000000000000000"; 
       x_416_tb <= "0000000000000000"; 
       x_417_tb <= "0000000000000000"; 
       x_418_tb <= "0000000000000000"; 
       x_419_tb <= "0000000000000000"; 
       x_420_tb <= "0000000000000000"; 
       x_421_tb <= "0000000000000000"; 
       x_422_tb <= "0000000000000000"; 
       x_423_tb <= "0000000000000000"; 
       x_424_tb <= "0000000000000000"; 
       x_425_tb <= "0000000000000000"; 
       x_426_tb <= "0000000000000000"; 
       x_427_tb <= "0000000000000000"; 
       x_428_tb <= "0000000000000000"; 
       x_429_tb <= "0000000000000000"; 
       x_430_tb <= "0000000000000000"; 
       x_431_tb <= "0000000000000000"; 
       x_432_tb <= "0000000000000000"; 
       x_433_tb <= "0000000010010110"; 
       x_434_tb <= "0000000011111110"; 
       x_435_tb <= "0000000011110100"; 
       x_436_tb <= "0000000000000000"; 
       x_437_tb <= "0000000000000000"; 
       x_438_tb <= "0000000000000000"; 
       x_439_tb <= "0000000000000000"; 
       x_440_tb <= "0000000000000000"; 
       x_441_tb <= "0000000000000000"; 
       x_442_tb <= "0000000000000000"; 
       x_443_tb <= "0000000000000000"; 
       x_444_tb <= "0000000000000000"; 
       x_445_tb <= "0000000000000000"; 
       x_446_tb <= "0000000000000000"; 
       x_447_tb <= "0000000000000000"; 
       x_448_tb <= "0000000000000000"; 
       x_449_tb <= "0000000000000000"; 
       x_450_tb <= "0000000000000000"; 
       x_451_tb <= "0000000000000000"; 
       x_452_tb <= "0000000000000000"; 
       x_453_tb <= "0000000000000000"; 
       x_454_tb <= "0000000000000000"; 
       x_455_tb <= "0000000000000000"; 
       x_456_tb <= "0000000000000000"; 
       x_457_tb <= "0000000000000000"; 
       x_458_tb <= "0000000000000000"; 
       x_459_tb <= "0000000000000000"; 
       x_460_tb <= "0000000000000000"; 
       x_461_tb <= "0000000011000100"; 
       x_462_tb <= "0000000011111110"; 
       x_463_tb <= "0000000010100101"; 
       x_464_tb <= "0000000000000000"; 
       x_465_tb <= "0000000000000000"; 
       x_466_tb <= "0000000000000000"; 
       x_467_tb <= "0000000000000000"; 
       x_468_tb <= "0000000000000000"; 
       x_469_tb <= "0000000000000000"; 
       x_470_tb <= "0000000000000000"; 
       x_471_tb <= "0000000000000000"; 
       x_472_tb <= "0000000000000000"; 
       x_473_tb <= "0000000000000000"; 
       x_474_tb <= "0000000000000000"; 
       x_475_tb <= "0000000000000000"; 
       x_476_tb <= "0000000000000000"; 
       x_477_tb <= "0000000000000000"; 
       x_478_tb <= "0000000000000000"; 
       x_479_tb <= "0000000000000000"; 
       x_480_tb <= "0000000000000000"; 
       x_481_tb <= "0000000000000000"; 
       x_482_tb <= "0000000000000000"; 
       x_483_tb <= "0000000000000000"; 
       x_484_tb <= "0000000000000000"; 
       x_485_tb <= "0000000000000000"; 
       x_486_tb <= "0000000000000000"; 
       x_487_tb <= "0000000000000000"; 
       x_488_tb <= "0000000000000000"; 
       x_489_tb <= "0000000010100110"; 
       x_490_tb <= "0000000011111110"; 
       x_491_tb <= "0000000011101001"; 
       x_492_tb <= "0000000000000000"; 
       x_493_tb <= "0000000000000000"; 
       x_494_tb <= "0000000000000000"; 
       x_495_tb <= "0000000000000000"; 
       x_496_tb <= "0000000000000000"; 
       x_497_tb <= "0000000000000000"; 
       x_498_tb <= "0000000000000000"; 
       x_499_tb <= "0000000000000000"; 
       x_500_tb <= "0000000000000000"; 
       x_501_tb <= "0000000000000000"; 
       x_502_tb <= "0000000000000000"; 
       x_503_tb <= "0000000000000000"; 
       x_504_tb <= "0000000000000000"; 
       x_505_tb <= "0000000000000000"; 
       x_506_tb <= "0000000000000000"; 
       x_507_tb <= "0000000000000000"; 
       x_508_tb <= "0000000000000000"; 
       x_509_tb <= "0000000000000000"; 
       x_510_tb <= "0000000000000000"; 
       x_511_tb <= "0000000000000000"; 
       x_512_tb <= "0000000000000000"; 
       x_513_tb <= "0000000000000000"; 
       x_514_tb <= "0000000000000000"; 
       x_515_tb <= "0000000000000000"; 
       x_516_tb <= "0000000000000000"; 
       x_517_tb <= "0000000000000000"; 
       x_518_tb <= "0000000011111110"; 
       x_519_tb <= "0000000011101001"; 
       x_520_tb <= "0000000000000000"; 
       x_521_tb <= "0000000000000000"; 
       x_522_tb <= "0000000000000000"; 
       x_523_tb <= "0000000000000000"; 
       x_524_tb <= "0000000000000000"; 
       x_525_tb <= "0000000000000000"; 
       x_526_tb <= "0000000000000000"; 
       x_527_tb <= "0000000000000000"; 
       x_528_tb <= "0000000000000000"; 
       x_529_tb <= "0000000000000000"; 
       x_530_tb <= "0000000000000000"; 
       x_531_tb <= "0000000000000000"; 
       x_532_tb <= "0000000000000000"; 
       x_533_tb <= "0000000000000000"; 
       x_534_tb <= "0000000000000000"; 
       x_535_tb <= "0000000000000000"; 
       x_536_tb <= "0000000000000000"; 
       x_537_tb <= "0000000000000000"; 
       x_538_tb <= "0000000000000000"; 
       x_539_tb <= "0000000000000000"; 
       x_540_tb <= "0000000000000000"; 
       x_541_tb <= "0000000000000000"; 
       x_542_tb <= "0000000000000000"; 
       x_543_tb <= "0000000000000000"; 
       x_544_tb <= "0000000000000000"; 
       x_545_tb <= "0000000000000000"; 
       x_546_tb <= "0000000011111111"; 
       x_547_tb <= "0000000011111110"; 
       x_548_tb <= "0000000010011100"; 
       x_549_tb <= "0000000000000000"; 
       x_550_tb <= "0000000000000000"; 
       x_551_tb <= "0000000000000000"; 
       x_552_tb <= "0000000000000000"; 
       x_553_tb <= "0000000000000000"; 
       x_554_tb <= "0000000000000000"; 
       x_555_tb <= "0000000000000000"; 
       x_556_tb <= "0000000000000000"; 
       x_557_tb <= "0000000000000000"; 
       x_558_tb <= "0000000000000000"; 
       x_559_tb <= "0000000000000000"; 
       x_560_tb <= "0000000000000000"; 
       x_561_tb <= "0000000000000000"; 
       x_562_tb <= "0000000000000000"; 
       x_563_tb <= "0000000000000000"; 
       x_564_tb <= "0000000000000000"; 
       x_565_tb <= "0000000000000000"; 
       x_566_tb <= "0000000000000000"; 
       x_567_tb <= "0000000000000000"; 
       x_568_tb <= "0000000000000000"; 
       x_569_tb <= "0000000000000000"; 
       x_570_tb <= "0000000000000000"; 
       x_571_tb <= "0000000000000000"; 
       x_572_tb <= "0000000000000000"; 
       x_573_tb <= "0000000000000000"; 
       x_574_tb <= "0000000011111110"; 
       x_575_tb <= "0000000011111101"; 
       x_576_tb <= "0000000010011100"; 
       x_577_tb <= "0000000000000000"; 
       x_578_tb <= "0000000000000000"; 
       x_579_tb <= "0000000000000000"; 
       x_580_tb <= "0000000000000000"; 
       x_581_tb <= "0000000000000000"; 
       x_582_tb <= "0000000000000000"; 
       x_583_tb <= "0000000000000000"; 
       x_584_tb <= "0000000000000000"; 
       x_585_tb <= "0000000000000000"; 
       x_586_tb <= "0000000000000000"; 
       x_587_tb <= "0000000000000000"; 
       x_588_tb <= "0000000000000000"; 
       x_589_tb <= "0000000000000000"; 
       x_590_tb <= "0000000000000000"; 
       x_591_tb <= "0000000000000000"; 
       x_592_tb <= "0000000000000000"; 
       x_593_tb <= "0000000000000000"; 
       x_594_tb <= "0000000000000000"; 
       x_595_tb <= "0000000000000000"; 
       x_596_tb <= "0000000000000000"; 
       x_597_tb <= "0000000000000000"; 
       x_598_tb <= "0000000000000000"; 
       x_599_tb <= "0000000000000000"; 
       x_600_tb <= "0000000000000000"; 
       x_601_tb <= "0000000000000000"; 
       x_602_tb <= "0000000011111110"; 
       x_603_tb <= "0000000011111101"; 
       x_604_tb <= "0000000010011100"; 
       x_605_tb <= "0000000000000000"; 
       x_606_tb <= "0000000000000000"; 
       x_607_tb <= "0000000000000000"; 
       x_608_tb <= "0000000000000000"; 
       x_609_tb <= "0000000000000000"; 
       x_610_tb <= "0000000000000000"; 
       x_611_tb <= "0000000000000000"; 
       x_612_tb <= "0000000000000000"; 
       x_613_tb <= "0000000000000000"; 
       x_614_tb <= "0000000000000000"; 
       x_615_tb <= "0000000000000000"; 
       x_616_tb <= "0000000000000000"; 
       x_617_tb <= "0000000000000000"; 
       x_618_tb <= "0000000000000000"; 
       x_619_tb <= "0000000000000000"; 
       x_620_tb <= "0000000000000000"; 
       x_621_tb <= "0000000000000000"; 
       x_622_tb <= "0000000000000000"; 
       x_623_tb <= "0000000000000000"; 
       x_624_tb <= "0000000000000000"; 
       x_625_tb <= "0000000000000000"; 
       x_626_tb <= "0000000000000000"; 
       x_627_tb <= "0000000000000000"; 
       x_628_tb <= "0000000000000000"; 
       x_629_tb <= "0000000000000000"; 
       x_630_tb <= "0000000011101110"; 
       x_631_tb <= "0000000011111101"; 
       x_632_tb <= "0000000010011100"; 
       x_633_tb <= "0000000000000000"; 
       x_634_tb <= "0000000000000000"; 
       x_635_tb <= "0000000000000000"; 
       x_636_tb <= "0000000000000000"; 
       x_637_tb <= "0000000000000000"; 
       x_638_tb <= "0000000000000000"; 
       x_639_tb <= "0000000000000000"; 
       x_640_tb <= "0000000000000000"; 
       x_641_tb <= "0000000000000000"; 
       x_642_tb <= "0000000000000000"; 
       x_643_tb <= "0000000000000000"; 
       x_644_tb <= "0000000000000000"; 
       x_645_tb <= "0000000000000000"; 
       x_646_tb <= "0000000000000000"; 
       x_647_tb <= "0000000000000000"; 
       x_648_tb <= "0000000000000000"; 
       x_649_tb <= "0000000000000000"; 
       x_650_tb <= "0000000000000000"; 
       x_651_tb <= "0000000000000000"; 
       x_652_tb <= "0000000000000000"; 
       x_653_tb <= "0000000000000000"; 
       x_654_tb <= "0000000000000000"; 
       x_655_tb <= "0000000000000000"; 
       x_656_tb <= "0000000000000000"; 
       x_657_tb <= "0000000000000000"; 
       x_658_tb <= "0000000010100010"; 
       x_659_tb <= "0000000011101101"; 
       x_660_tb <= "0000000010010000"; 
       x_661_tb <= "0000000000000000"; 
       x_662_tb <= "0000000000000000"; 
       x_663_tb <= "0000000000000000"; 
       x_664_tb <= "0000000000000000"; 
       x_665_tb <= "0000000000000000"; 
       x_666_tb <= "0000000000000000"; 
       x_667_tb <= "0000000000000000"; 
       x_668_tb <= "0000000000000000"; 
       x_669_tb <= "0000000000000000"; 
       x_670_tb <= "0000000000000000"; 
       x_671_tb <= "0000000000000000"; 
       x_672_tb <= "0000000000000000"; 
       x_673_tb <= "0000000000000000"; 
       x_674_tb <= "0000000000000000"; 
       x_675_tb <= "0000000000000000"; 
       x_676_tb <= "0000000000000000"; 
       x_677_tb <= "0000000000000000"; 
       x_678_tb <= "0000000000000000"; 
       x_679_tb <= "0000000000000000"; 
       x_680_tb <= "0000000000000000"; 
       x_681_tb <= "0000000000000000"; 
       x_682_tb <= "0000000000000000"; 
       x_683_tb <= "0000000000000000"; 
       x_684_tb <= "0000000000000000"; 
       x_685_tb <= "0000000000000000"; 
       x_686_tb <= "0000000000000000"; 
       x_687_tb <= "0000000000000000"; 
       x_688_tb <= "0000000000000000"; 
       x_689_tb <= "0000000000000000"; 
       x_690_tb <= "0000000000000000"; 
       x_691_tb <= "0000000000000000"; 
       x_692_tb <= "0000000000000000"; 
       x_693_tb <= "0000000000000000"; 
       x_694_tb <= "0000000000000000"; 
       x_695_tb <= "0000000000000000"; 
       x_696_tb <= "0000000000000000"; 
       x_697_tb <= "0000000000000000"; 
       x_698_tb <= "0000000000000000"; 
       x_699_tb <= "0000000000000000"; 
       x_700_tb <= "0000000000000000"; 
       x_701_tb <= "0000000000000000"; 
       x_702_tb <= "0000000000000000"; 
       x_703_tb <= "0000000000000000"; 
       x_704_tb <= "0000000000000000"; 
       x_705_tb <= "0000000000000000"; 
       x_706_tb <= "0000000000000000"; 
       x_707_tb <= "0000000000000000"; 
       x_708_tb <= "0000000000000000"; 
       x_709_tb <= "0000000000000000"; 
       x_710_tb <= "0000000000000000"; 
       x_711_tb <= "0000000000000000"; 
       x_712_tb <= "0000000000000000"; 
       x_713_tb <= "0000000000000000"; 
       x_714_tb <= "0000000000000000"; 
       x_715_tb <= "0000000000000000"; 
       x_716_tb <= "0000000000000000"; 
       x_717_tb <= "0000000000000000"; 
       x_718_tb <= "0000000000000000"; 
       x_719_tb <= "0000000000000000"; 
       x_720_tb <= "0000000000000000"; 
       x_721_tb <= "0000000000000000"; 
       x_722_tb <= "0000000000000000"; 
       x_723_tb <= "0000000000000000"; 
       x_724_tb <= "0000000000000000"; 
       x_725_tb <= "0000000000000000"; 
       x_726_tb <= "0000000000000000"; 
       x_727_tb <= "0000000000000000"; 
       x_728_tb <= "0000000000000000"; 
       x_729_tb <= "0000000000000000"; 
       x_730_tb <= "0000000000000000"; 
       x_731_tb <= "0000000000000000"; 
       x_732_tb <= "0000000000000000"; 
       x_733_tb <= "0000000000000000"; 
       x_734_tb <= "0000000000000000"; 
       x_735_tb <= "0000000000000000"; 
       x_736_tb <= "0000000000000000"; 
       x_737_tb <= "0000000000000000"; 
       x_738_tb <= "0000000000000000"; 
       x_739_tb <= "0000000000000000"; 
       x_740_tb <= "0000000000000000"; 
       x_741_tb <= "0000000000000000"; 
       x_742_tb <= "0000000000000000"; 
       x_743_tb <= "0000000000000000"; 
       x_744_tb <= "0000000000000000"; 
       x_745_tb <= "0000000000000000"; 
       x_746_tb <= "0000000000000000"; 
       x_747_tb <= "0000000000000000"; 
       x_748_tb <= "0000000000000000"; 
       x_749_tb <= "0000000000000000"; 
       x_750_tb <= "0000000000000000"; 
       x_751_tb <= "0000000000000000"; 
       x_752_tb <= "0000000000000000"; 
       x_753_tb <= "0000000000000000"; 
       x_754_tb <= "0000000000000000"; 
       x_755_tb <= "0000000000000000"; 
       x_756_tb <= "0000000000000000"; 
       x_757_tb <= "0000000000000000"; 
       x_758_tb <= "0000000000000000"; 
       x_759_tb <= "0000000000000000"; 
       x_760_tb <= "0000000000000000"; 
       x_761_tb <= "0000000000000000"; 
       x_762_tb <= "0000000000000000"; 
       x_763_tb <= "0000000000000000"; 
       x_764_tb <= "0000000000000000"; 
       x_765_tb <= "0000000000000000"; 
       x_766_tb <= "0000000000000000"; 
       x_767_tb <= "0000000000000000"; 
       x_768_tb <= "0000000000000000"; 
       x_769_tb <= "0000000000000000"; 
       x_770_tb <= "0000000000000000"; 
       x_771_tb <= "0000000000000000"; 
       x_772_tb <= "0000000000000000"; 
       x_773_tb <= "0000000000000000"; 
       x_774_tb <= "0000000000000000"; 
       x_775_tb <= "0000000000000000"; 
       x_776_tb <= "0000000000000000"; 
       x_777_tb <= "0000000000000000"; 
       x_778_tb <= "0000000000000000"; 
       x_779_tb <= "0000000000000000"; 
       x_780_tb <= "0000000000000000"; 
       x_781_tb <= "0000000000000000"; 
       x_782_tb <= "0000000000000000"; 
       x_783_tb <= "0000000000000000"; 
    wait for 750 ns;
   wait ;
    end process ;
end Behavioral ;
