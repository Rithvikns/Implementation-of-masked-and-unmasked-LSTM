library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity lstm_layer is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_0 : out STD_LOGIC_VECTOR(15 downto 0);
        y_1 : out STD_LOGIC_VECTOR(15 downto 0);
        y_2 : out STD_LOGIC_VECTOR(15 downto 0);
        y_3 : out STD_LOGIC_VECTOR(15 downto 0);
        y_4 : out STD_LOGIC_VECTOR(15 downto 0);
        y_5 : out STD_LOGIC_VECTOR(15 downto 0);
        y_6 : out STD_LOGIC_VECTOR(15 downto 0);
        y_7 : out STD_LOGIC_VECTOR(15 downto 0);
        y_8 : out STD_LOGIC_VECTOR(15 downto 0);
        y_9 : out STD_LOGIC_VECTOR(15 downto 0);
        y_10 : out STD_LOGIC_VECTOR(15 downto 0);
        y_11 : out STD_LOGIC_VECTOR(15 downto 0);
        y_12 : out STD_LOGIC_VECTOR(15 downto 0);
        y_13 : out STD_LOGIC_VECTOR(15 downto 0);
        y_14 : out STD_LOGIC_VECTOR(15 downto 0);
        y_15 : out STD_LOGIC_VECTOR(15 downto 0);
        y_16 : out STD_LOGIC_VECTOR(15 downto 0);
        y_17 : out STD_LOGIC_VECTOR(15 downto 0);
        y_18 : out STD_LOGIC_VECTOR(15 downto 0);
        y_19 : out STD_LOGIC_VECTOR(15 downto 0);
        y_20 : out STD_LOGIC_VECTOR(15 downto 0);
        y_21 : out STD_LOGIC_VECTOR(15 downto 0);
        y_22 : out STD_LOGIC_VECTOR(15 downto 0);
        y_23 : out STD_LOGIC_VECTOR(15 downto 0);
        y_24 : out STD_LOGIC_VECTOR(15 downto 0);
        y_25 : out STD_LOGIC_VECTOR(15 downto 0);
        y_26 : out STD_LOGIC_VECTOR(15 downto 0);
        y_27 : out STD_LOGIC_VECTOR(15 downto 0);
        y_28 : out STD_LOGIC_VECTOR(15 downto 0);
        y_29 : out STD_LOGIC_VECTOR(15 downto 0);
        y_30 : out STD_LOGIC_VECTOR(15 downto 0);
        y_31 : out STD_LOGIC_VECTOR(15 downto 0);
        y_32 : out STD_LOGIC_VECTOR(15 downto 0);
        y_33 : out STD_LOGIC_VECTOR(15 downto 0);
        y_34 : out STD_LOGIC_VECTOR(15 downto 0);
        y_35 : out STD_LOGIC_VECTOR(15 downto 0);
        y_36 : out STD_LOGIC_VECTOR(15 downto 0);
        y_37 : out STD_LOGIC_VECTOR(15 downto 0);
        y_38 : out STD_LOGIC_VECTOR(15 downto 0);
        y_39 : out STD_LOGIC_VECTOR(15 downto 0);
        y_40 : out STD_LOGIC_VECTOR(15 downto 0);
        y_41 : out STD_LOGIC_VECTOR(15 downto 0);
        y_42 : out STD_LOGIC_VECTOR(15 downto 0);
        y_43 : out STD_LOGIC_VECTOR(15 downto 0);
        y_44 : out STD_LOGIC_VECTOR(15 downto 0);
        y_45 : out STD_LOGIC_VECTOR(15 downto 0);
        y_46 : out STD_LOGIC_VECTOR(15 downto 0);
        y_47 : out STD_LOGIC_VECTOR(15 downto 0);
        y_48 : out STD_LOGIC_VECTOR(15 downto 0);
        y_49 : out STD_LOGIC_VECTOR(15 downto 0);
        y_50 : out STD_LOGIC_VECTOR(15 downto 0);
        y_51 : out STD_LOGIC_VECTOR(15 downto 0);
        y_52 : out STD_LOGIC_VECTOR(15 downto 0);
        y_53 : out STD_LOGIC_VECTOR(15 downto 0);
        y_54 : out STD_LOGIC_VECTOR(15 downto 0);
        y_55 : out STD_LOGIC_VECTOR(15 downto 0);
        y_56 : out STD_LOGIC_VECTOR(15 downto 0);
        y_57 : out STD_LOGIC_VECTOR(15 downto 0);
        y_58 : out STD_LOGIC_VECTOR(15 downto 0);
        y_59 : out STD_LOGIC_VECTOR(15 downto 0);
        y_60 : out STD_LOGIC_VECTOR(15 downto 0);
        y_61 : out STD_LOGIC_VECTOR(15 downto 0);
        y_62 : out STD_LOGIC_VECTOR(15 downto 0);
        y_63 : out STD_LOGIC_VECTOR(15 downto 0);
        y_64 : out STD_LOGIC_VECTOR(15 downto 0);
        y_65 : out STD_LOGIC_VECTOR(15 downto 0);
        y_66 : out STD_LOGIC_VECTOR(15 downto 0);
        y_67 : out STD_LOGIC_VECTOR(15 downto 0);
        y_68 : out STD_LOGIC_VECTOR(15 downto 0);
        y_69 : out STD_LOGIC_VECTOR(15 downto 0);
        y_70 : out STD_LOGIC_VECTOR(15 downto 0);
        y_71 : out STD_LOGIC_VECTOR(15 downto 0);
        y_72 : out STD_LOGIC_VECTOR(15 downto 0);
        y_73 : out STD_LOGIC_VECTOR(15 downto 0);
        y_74 : out STD_LOGIC_VECTOR(15 downto 0);
        y_75 : out STD_LOGIC_VECTOR(15 downto 0);
        y_76 : out STD_LOGIC_VECTOR(15 downto 0);
        y_77 : out STD_LOGIC_VECTOR(15 downto 0);
        y_78 : out STD_LOGIC_VECTOR(15 downto 0);
        y_79 : out STD_LOGIC_VECTOR(15 downto 0);
        y_80 : out STD_LOGIC_VECTOR(15 downto 0);
        y_81 : out STD_LOGIC_VECTOR(15 downto 0);
        y_82 : out STD_LOGIC_VECTOR(15 downto 0);
        y_83 : out STD_LOGIC_VECTOR(15 downto 0);
        y_84 : out STD_LOGIC_VECTOR(15 downto 0);
        y_85 : out STD_LOGIC_VECTOR(15 downto 0);
        y_86 : out STD_LOGIC_VECTOR(15 downto 0);
        y_87 : out STD_LOGIC_VECTOR(15 downto 0);
        y_88 : out STD_LOGIC_VECTOR(15 downto 0);
        y_89 : out STD_LOGIC_VECTOR(15 downto 0);
        y_90 : out STD_LOGIC_VECTOR(15 downto 0);
        y_91 : out STD_LOGIC_VECTOR(15 downto 0);
        y_92 : out STD_LOGIC_VECTOR(15 downto 0);
        y_93 : out STD_LOGIC_VECTOR(15 downto 0);
        y_94 : out STD_LOGIC_VECTOR(15 downto 0);
        y_95 : out STD_LOGIC_VECTOR(15 downto 0);
        y_96 : out STD_LOGIC_VECTOR(15 downto 0);
        y_97 : out STD_LOGIC_VECTOR(15 downto 0);
        y_98 : out STD_LOGIC_VECTOR(15 downto 0);
        y_99 : out STD_LOGIC_VECTOR(15 downto 0);
        y_100 : out STD_LOGIC_VECTOR(15 downto 0);
        y_101 : out STD_LOGIC_VECTOR(15 downto 0);
        y_102 : out STD_LOGIC_VECTOR(15 downto 0);
        y_103 : out STD_LOGIC_VECTOR(15 downto 0);
        y_104 : out STD_LOGIC_VECTOR(15 downto 0);
        y_105 : out STD_LOGIC_VECTOR(15 downto 0);
        y_106 : out STD_LOGIC_VECTOR(15 downto 0);
        y_107 : out STD_LOGIC_VECTOR(15 downto 0);
        y_108 : out STD_LOGIC_VECTOR(15 downto 0);
        y_109 : out STD_LOGIC_VECTOR(15 downto 0);
        y_110 : out STD_LOGIC_VECTOR(15 downto 0);
        y_111 : out STD_LOGIC_VECTOR(15 downto 0);
        y_112 : out STD_LOGIC_VECTOR(15 downto 0);
        y_113 : out STD_LOGIC_VECTOR(15 downto 0);
        y_114 : out STD_LOGIC_VECTOR(15 downto 0);
        y_115 : out STD_LOGIC_VECTOR(15 downto 0);
        y_116 : out STD_LOGIC_VECTOR(15 downto 0);
        y_117 : out STD_LOGIC_VECTOR(15 downto 0);
        y_118 : out STD_LOGIC_VECTOR(15 downto 0);
        y_119 : out STD_LOGIC_VECTOR(15 downto 0);
        y_120 : out STD_LOGIC_VECTOR(15 downto 0);
        y_121 : out STD_LOGIC_VECTOR(15 downto 0);
        y_122 : out STD_LOGIC_VECTOR(15 downto 0);
        y_123 : out STD_LOGIC_VECTOR(15 downto 0);
        y_124 : out STD_LOGIC_VECTOR(15 downto 0);
        y_125 : out STD_LOGIC_VECTOR(15 downto 0);
        y_126 : out STD_LOGIC_VECTOR(15 downto 0);
        y_127 : out STD_LOGIC_VECTOR(15 downto 0);
        y_128 : out STD_LOGIC_VECTOR(15 downto 0);
        y_129 : out STD_LOGIC_VECTOR(15 downto 0);
        y_130 : out STD_LOGIC_VECTOR(15 downto 0);
        y_131 : out STD_LOGIC_VECTOR(15 downto 0);
        y_132 : out STD_LOGIC_VECTOR(15 downto 0);
        y_133 : out STD_LOGIC_VECTOR(15 downto 0);
        y_134 : out STD_LOGIC_VECTOR(15 downto 0);
        y_135 : out STD_LOGIC_VECTOR(15 downto 0);
        y_136 : out STD_LOGIC_VECTOR(15 downto 0);
        y_137 : out STD_LOGIC_VECTOR(15 downto 0);
        y_138 : out STD_LOGIC_VECTOR(15 downto 0);
        y_139 : out STD_LOGIC_VECTOR(15 downto 0);
        y_140 : out STD_LOGIC_VECTOR(15 downto 0);
        y_141 : out STD_LOGIC_VECTOR(15 downto 0);
        y_142 : out STD_LOGIC_VECTOR(15 downto 0);
        y_143 : out STD_LOGIC_VECTOR(15 downto 0);
        y_144 : out STD_LOGIC_VECTOR(15 downto 0);
        y_145 : out STD_LOGIC_VECTOR(15 downto 0);
        y_146 : out STD_LOGIC_VECTOR(15 downto 0);
        y_147 : out STD_LOGIC_VECTOR(15 downto 0);
        y_148 : out STD_LOGIC_VECTOR(15 downto 0);
        y_149 : out STD_LOGIC_VECTOR(15 downto 0);
        y_150 : out STD_LOGIC_VECTOR(15 downto 0);
        y_151 : out STD_LOGIC_VECTOR(15 downto 0);
        y_152 : out STD_LOGIC_VECTOR(15 downto 0);
        y_153 : out STD_LOGIC_VECTOR(15 downto 0);
        y_154 : out STD_LOGIC_VECTOR(15 downto 0);
        y_155 : out STD_LOGIC_VECTOR(15 downto 0);
        y_156 : out STD_LOGIC_VECTOR(15 downto 0);
        y_157 : out STD_LOGIC_VECTOR(15 downto 0);
        y_158 : out STD_LOGIC_VECTOR(15 downto 0);
        y_159 : out STD_LOGIC_VECTOR(15 downto 0);
        y_160 : out STD_LOGIC_VECTOR(15 downto 0);
        y_161 : out STD_LOGIC_VECTOR(15 downto 0);
        y_162 : out STD_LOGIC_VECTOR(15 downto 0);
        y_163 : out STD_LOGIC_VECTOR(15 downto 0);
        y_164 : out STD_LOGIC_VECTOR(15 downto 0);
        y_165 : out STD_LOGIC_VECTOR(15 downto 0);
        y_166 : out STD_LOGIC_VECTOR(15 downto 0);
        y_167 : out STD_LOGIC_VECTOR(15 downto 0);
        y_168 : out STD_LOGIC_VECTOR(15 downto 0);
        y_169 : out STD_LOGIC_VECTOR(15 downto 0);
        y_170 : out STD_LOGIC_VECTOR(15 downto 0);
        y_171 : out STD_LOGIC_VECTOR(15 downto 0);
        y_172 : out STD_LOGIC_VECTOR(15 downto 0);
        y_173 : out STD_LOGIC_VECTOR(15 downto 0);
        y_174 : out STD_LOGIC_VECTOR(15 downto 0);
        y_175 : out STD_LOGIC_VECTOR(15 downto 0);
        y_176 : out STD_LOGIC_VECTOR(15 downto 0);
        y_177 : out STD_LOGIC_VECTOR(15 downto 0);
        y_178 : out STD_LOGIC_VECTOR(15 downto 0);
        y_179 : out STD_LOGIC_VECTOR(15 downto 0);
        y_180 : out STD_LOGIC_VECTOR(15 downto 0);
        y_181 : out STD_LOGIC_VECTOR(15 downto 0);
        y_182 : out STD_LOGIC_VECTOR(15 downto 0);
        y_183 : out STD_LOGIC_VECTOR(15 downto 0);
        y_184 : out STD_LOGIC_VECTOR(15 downto 0);
        y_185 : out STD_LOGIC_VECTOR(15 downto 0);
        y_186 : out STD_LOGIC_VECTOR(15 downto 0);
        y_187 : out STD_LOGIC_VECTOR(15 downto 0);
        y_188 : out STD_LOGIC_VECTOR(15 downto 0);
        y_189 : out STD_LOGIC_VECTOR(15 downto 0);
        y_190 : out STD_LOGIC_VECTOR(15 downto 0);
        y_191 : out STD_LOGIC_VECTOR(15 downto 0);
        y_192 : out STD_LOGIC_VECTOR(15 downto 0);
        y_193 : out STD_LOGIC_VECTOR(15 downto 0);
        y_194 : out STD_LOGIC_VECTOR(15 downto 0);
        y_195 : out STD_LOGIC_VECTOR(15 downto 0);
        y_196 : out STD_LOGIC_VECTOR(15 downto 0);
        y_197 : out STD_LOGIC_VECTOR(15 downto 0);
        y_198 : out STD_LOGIC_VECTOR(15 downto 0);
        y_199 : out STD_LOGIC_VECTOR(15 downto 0);
        y_200 : out STD_LOGIC_VECTOR(15 downto 0);
        y_201 : out STD_LOGIC_VECTOR(15 downto 0);
        y_202 : out STD_LOGIC_VECTOR(15 downto 0);
        y_203 : out STD_LOGIC_VECTOR(15 downto 0);
        y_204 : out STD_LOGIC_VECTOR(15 downto 0);
        y_205 : out STD_LOGIC_VECTOR(15 downto 0);
        y_206 : out STD_LOGIC_VECTOR(15 downto 0);
        y_207 : out STD_LOGIC_VECTOR(15 downto 0);
        y_208 : out STD_LOGIC_VECTOR(15 downto 0);
        y_209 : out STD_LOGIC_VECTOR(15 downto 0);
        y_210 : out STD_LOGIC_VECTOR(15 downto 0);
        y_211 : out STD_LOGIC_VECTOR(15 downto 0);
        y_212 : out STD_LOGIC_VECTOR(15 downto 0);
        y_213 : out STD_LOGIC_VECTOR(15 downto 0);
        y_214 : out STD_LOGIC_VECTOR(15 downto 0);
        y_215 : out STD_LOGIC_VECTOR(15 downto 0);
        y_216 : out STD_LOGIC_VECTOR(15 downto 0);
        y_217 : out STD_LOGIC_VECTOR(15 downto 0);
        y_218 : out STD_LOGIC_VECTOR(15 downto 0);
        y_219 : out STD_LOGIC_VECTOR(15 downto 0);
        y_220 : out STD_LOGIC_VECTOR(15 downto 0);
        y_221 : out STD_LOGIC_VECTOR(15 downto 0);
        y_222 : out STD_LOGIC_VECTOR(15 downto 0);
        y_223 : out STD_LOGIC_VECTOR(15 downto 0);
        y_224 : out STD_LOGIC_VECTOR(15 downto 0);
        y_225 : out STD_LOGIC_VECTOR(15 downto 0);
        y_226 : out STD_LOGIC_VECTOR(15 downto 0);
        y_227 : out STD_LOGIC_VECTOR(15 downto 0);
        y_228 : out STD_LOGIC_VECTOR(15 downto 0);
        y_229 : out STD_LOGIC_VECTOR(15 downto 0);
        y_230 : out STD_LOGIC_VECTOR(15 downto 0);
        y_231 : out STD_LOGIC_VECTOR(15 downto 0);
        y_232 : out STD_LOGIC_VECTOR(15 downto 0);
        y_233 : out STD_LOGIC_VECTOR(15 downto 0);
        y_234 : out STD_LOGIC_VECTOR(15 downto 0);
        y_235 : out STD_LOGIC_VECTOR(15 downto 0);
        y_236 : out STD_LOGIC_VECTOR(15 downto 0);
        y_237 : out STD_LOGIC_VECTOR(15 downto 0);
        y_238 : out STD_LOGIC_VECTOR(15 downto 0);
        y_239 : out STD_LOGIC_VECTOR(15 downto 0);
        y_240 : out STD_LOGIC_VECTOR(15 downto 0);
        y_241 : out STD_LOGIC_VECTOR(15 downto 0);
        y_242 : out STD_LOGIC_VECTOR(15 downto 0);
        y_243 : out STD_LOGIC_VECTOR(15 downto 0);
        y_244 : out STD_LOGIC_VECTOR(15 downto 0);
        y_245 : out STD_LOGIC_VECTOR(15 downto 0);
        y_246 : out STD_LOGIC_VECTOR(15 downto 0);
        y_247 : out STD_LOGIC_VECTOR(15 downto 0);
        y_248 : out STD_LOGIC_VECTOR(15 downto 0);
        y_249 : out STD_LOGIC_VECTOR(15 downto 0);
        y_250 : out STD_LOGIC_VECTOR(15 downto 0);
        y_251 : out STD_LOGIC_VECTOR(15 downto 0);
        y_252 : out STD_LOGIC_VECTOR(15 downto 0);
        y_253 : out STD_LOGIC_VECTOR(15 downto 0);
        y_254 : out STD_LOGIC_VECTOR(15 downto 0);
        y_255 : out STD_LOGIC_VECTOR(15 downto 0);
        y_256 : out STD_LOGIC_VECTOR(15 downto 0);
        y_257 : out STD_LOGIC_VECTOR(15 downto 0);
        y_258 : out STD_LOGIC_VECTOR(15 downto 0);
        y_259 : out STD_LOGIC_VECTOR(15 downto 0);
        y_260 : out STD_LOGIC_VECTOR(15 downto 0);
        y_261 : out STD_LOGIC_VECTOR(15 downto 0);
        y_262 : out STD_LOGIC_VECTOR(15 downto 0);
        y_263 : out STD_LOGIC_VECTOR(15 downto 0);
        y_264 : out STD_LOGIC_VECTOR(15 downto 0);
        y_265 : out STD_LOGIC_VECTOR(15 downto 0);
        y_266 : out STD_LOGIC_VECTOR(15 downto 0);
        y_267 : out STD_LOGIC_VECTOR(15 downto 0);
        y_268 : out STD_LOGIC_VECTOR(15 downto 0);
        y_269 : out STD_LOGIC_VECTOR(15 downto 0);
        y_270 : out STD_LOGIC_VECTOR(15 downto 0);
        y_271 : out STD_LOGIC_VECTOR(15 downto 0);
        y_272 : out STD_LOGIC_VECTOR(15 downto 0);
        y_273 : out STD_LOGIC_VECTOR(15 downto 0);
        y_274 : out STD_LOGIC_VECTOR(15 downto 0);
        y_275 : out STD_LOGIC_VECTOR(15 downto 0);
        y_276 : out STD_LOGIC_VECTOR(15 downto 0);
        y_277 : out STD_LOGIC_VECTOR(15 downto 0);
        y_278 : out STD_LOGIC_VECTOR(15 downto 0);
        y_279 : out STD_LOGIC_VECTOR(15 downto 0);
        y_280 : out STD_LOGIC_VECTOR(15 downto 0);
        y_281 : out STD_LOGIC_VECTOR(15 downto 0);
        y_282 : out STD_LOGIC_VECTOR(15 downto 0);
        y_283 : out STD_LOGIC_VECTOR(15 downto 0);
        y_284 : out STD_LOGIC_VECTOR(15 downto 0);
        y_285 : out STD_LOGIC_VECTOR(15 downto 0);
        y_286 : out STD_LOGIC_VECTOR(15 downto 0);
        y_287 : out STD_LOGIC_VECTOR(15 downto 0);
        y_288 : out STD_LOGIC_VECTOR(15 downto 0);
        y_289 : out STD_LOGIC_VECTOR(15 downto 0);
        y_290 : out STD_LOGIC_VECTOR(15 downto 0);
        y_291 : out STD_LOGIC_VECTOR(15 downto 0);
        y_292 : out STD_LOGIC_VECTOR(15 downto 0);
        y_293 : out STD_LOGIC_VECTOR(15 downto 0);
        y_294 : out STD_LOGIC_VECTOR(15 downto 0);
        y_295 : out STD_LOGIC_VECTOR(15 downto 0);
        y_296 : out STD_LOGIC_VECTOR(15 downto 0);
        y_297 : out STD_LOGIC_VECTOR(15 downto 0);
        y_298 : out STD_LOGIC_VECTOR(15 downto 0);
        y_299 : out STD_LOGIC_VECTOR(15 downto 0);
        y_300 : out STD_LOGIC_VECTOR(15 downto 0);
        y_301 : out STD_LOGIC_VECTOR(15 downto 0);
        y_302 : out STD_LOGIC_VECTOR(15 downto 0);
        y_303 : out STD_LOGIC_VECTOR(15 downto 0);
        y_304 : out STD_LOGIC_VECTOR(15 downto 0);
        y_305 : out STD_LOGIC_VECTOR(15 downto 0);
        y_306 : out STD_LOGIC_VECTOR(15 downto 0);
        y_307 : out STD_LOGIC_VECTOR(15 downto 0);
        y_308 : out STD_LOGIC_VECTOR(15 downto 0);
        y_309 : out STD_LOGIC_VECTOR(15 downto 0);
        y_310 : out STD_LOGIC_VECTOR(15 downto 0);
        y_311 : out STD_LOGIC_VECTOR(15 downto 0);
        y_312 : out STD_LOGIC_VECTOR(15 downto 0);
        y_313 : out STD_LOGIC_VECTOR(15 downto 0);
        y_314 : out STD_LOGIC_VECTOR(15 downto 0);
        y_315 : out STD_LOGIC_VECTOR(15 downto 0);
        y_316 : out STD_LOGIC_VECTOR(15 downto 0);
        y_317 : out STD_LOGIC_VECTOR(15 downto 0);
        y_318 : out STD_LOGIC_VECTOR(15 downto 0);
        y_319 : out STD_LOGIC_VECTOR(15 downto 0);
        y_320 : out STD_LOGIC_VECTOR(15 downto 0);
        y_321 : out STD_LOGIC_VECTOR(15 downto 0);
        y_322 : out STD_LOGIC_VECTOR(15 downto 0);
        y_323 : out STD_LOGIC_VECTOR(15 downto 0);
        y_324 : out STD_LOGIC_VECTOR(15 downto 0);
        y_325 : out STD_LOGIC_VECTOR(15 downto 0);
        y_326 : out STD_LOGIC_VECTOR(15 downto 0);
        y_327 : out STD_LOGIC_VECTOR(15 downto 0);
        y_328 : out STD_LOGIC_VECTOR(15 downto 0);
        y_329 : out STD_LOGIC_VECTOR(15 downto 0);
        y_330 : out STD_LOGIC_VECTOR(15 downto 0);
        y_331 : out STD_LOGIC_VECTOR(15 downto 0);
        y_332 : out STD_LOGIC_VECTOR(15 downto 0);
        y_333 : out STD_LOGIC_VECTOR(15 downto 0);
        y_334 : out STD_LOGIC_VECTOR(15 downto 0);
        y_335 : out STD_LOGIC_VECTOR(15 downto 0);
        y_336 : out STD_LOGIC_VECTOR(15 downto 0);
        y_337 : out STD_LOGIC_VECTOR(15 downto 0);
        y_338 : out STD_LOGIC_VECTOR(15 downto 0);
        y_339 : out STD_LOGIC_VECTOR(15 downto 0);
        y_340 : out STD_LOGIC_VECTOR(15 downto 0);
        y_341 : out STD_LOGIC_VECTOR(15 downto 0);
        y_342 : out STD_LOGIC_VECTOR(15 downto 0);
        y_343 : out STD_LOGIC_VECTOR(15 downto 0);
        y_344 : out STD_LOGIC_VECTOR(15 downto 0);
        y_345 : out STD_LOGIC_VECTOR(15 downto 0);
        y_346 : out STD_LOGIC_VECTOR(15 downto 0);
        y_347 : out STD_LOGIC_VECTOR(15 downto 0);
        y_348 : out STD_LOGIC_VECTOR(15 downto 0);
        y_349 : out STD_LOGIC_VECTOR(15 downto 0);
        y_350 : out STD_LOGIC_VECTOR(15 downto 0);
        y_351 : out STD_LOGIC_VECTOR(15 downto 0);
        y_352 : out STD_LOGIC_VECTOR(15 downto 0);
        y_353 : out STD_LOGIC_VECTOR(15 downto 0);
        y_354 : out STD_LOGIC_VECTOR(15 downto 0);
        y_355 : out STD_LOGIC_VECTOR(15 downto 0);
        y_356 : out STD_LOGIC_VECTOR(15 downto 0);
        y_357 : out STD_LOGIC_VECTOR(15 downto 0);
        y_358 : out STD_LOGIC_VECTOR(15 downto 0);
        y_359 : out STD_LOGIC_VECTOR(15 downto 0);
        y_360 : out STD_LOGIC_VECTOR(15 downto 0);
        y_361 : out STD_LOGIC_VECTOR(15 downto 0);
        y_362 : out STD_LOGIC_VECTOR(15 downto 0);
        y_363 : out STD_LOGIC_VECTOR(15 downto 0);
        y_364 : out STD_LOGIC_VECTOR(15 downto 0);
        y_365 : out STD_LOGIC_VECTOR(15 downto 0);
        y_366 : out STD_LOGIC_VECTOR(15 downto 0);
        y_367 : out STD_LOGIC_VECTOR(15 downto 0);
        y_368 : out STD_LOGIC_VECTOR(15 downto 0);
        y_369 : out STD_LOGIC_VECTOR(15 downto 0);
        y_370 : out STD_LOGIC_VECTOR(15 downto 0);
        y_371 : out STD_LOGIC_VECTOR(15 downto 0);
        y_372 : out STD_LOGIC_VECTOR(15 downto 0);
        y_373 : out STD_LOGIC_VECTOR(15 downto 0);
        y_374 : out STD_LOGIC_VECTOR(15 downto 0);
        y_375 : out STD_LOGIC_VECTOR(15 downto 0);
        y_376 : out STD_LOGIC_VECTOR(15 downto 0);
        y_377 : out STD_LOGIC_VECTOR(15 downto 0);
        y_378 : out STD_LOGIC_VECTOR(15 downto 0);
        y_379 : out STD_LOGIC_VECTOR(15 downto 0);
        y_380 : out STD_LOGIC_VECTOR(15 downto 0);
        y_381 : out STD_LOGIC_VECTOR(15 downto 0);
        y_382 : out STD_LOGIC_VECTOR(15 downto 0);
        y_383 : out STD_LOGIC_VECTOR(15 downto 0);
        y_384 : out STD_LOGIC_VECTOR(15 downto 0);
        y_385 : out STD_LOGIC_VECTOR(15 downto 0);
        y_386 : out STD_LOGIC_VECTOR(15 downto 0);
        y_387 : out STD_LOGIC_VECTOR(15 downto 0);
        y_388 : out STD_LOGIC_VECTOR(15 downto 0);
        y_389 : out STD_LOGIC_VECTOR(15 downto 0);
        y_390 : out STD_LOGIC_VECTOR(15 downto 0);
        y_391 : out STD_LOGIC_VECTOR(15 downto 0);
        y_392 : out STD_LOGIC_VECTOR(15 downto 0);
        y_393 : out STD_LOGIC_VECTOR(15 downto 0);
        y_394 : out STD_LOGIC_VECTOR(15 downto 0);
        y_395 : out STD_LOGIC_VECTOR(15 downto 0);
        y_396 : out STD_LOGIC_VECTOR(15 downto 0);
        y_397 : out STD_LOGIC_VECTOR(15 downto 0);
        y_398 : out STD_LOGIC_VECTOR(15 downto 0);
        y_399 : out STD_LOGIC_VECTOR(15 downto 0);
        y_400 : out STD_LOGIC_VECTOR(15 downto 0);
        y_401 : out STD_LOGIC_VECTOR(15 downto 0);
        y_402 : out STD_LOGIC_VECTOR(15 downto 0);
        y_403 : out STD_LOGIC_VECTOR(15 downto 0);
        y_404 : out STD_LOGIC_VECTOR(15 downto 0);
        y_405 : out STD_LOGIC_VECTOR(15 downto 0);
        y_406 : out STD_LOGIC_VECTOR(15 downto 0);
        y_407 : out STD_LOGIC_VECTOR(15 downto 0);
        y_408 : out STD_LOGIC_VECTOR(15 downto 0);
        y_409 : out STD_LOGIC_VECTOR(15 downto 0);
        y_410 : out STD_LOGIC_VECTOR(15 downto 0);
        y_411 : out STD_LOGIC_VECTOR(15 downto 0);
        y_412 : out STD_LOGIC_VECTOR(15 downto 0);
        y_413 : out STD_LOGIC_VECTOR(15 downto 0);
        y_414 : out STD_LOGIC_VECTOR(15 downto 0);
        y_415 : out STD_LOGIC_VECTOR(15 downto 0);
        y_416 : out STD_LOGIC_VECTOR(15 downto 0);
        y_417 : out STD_LOGIC_VECTOR(15 downto 0);
        y_418 : out STD_LOGIC_VECTOR(15 downto 0);
        y_419 : out STD_LOGIC_VECTOR(15 downto 0);
        y_420 : out STD_LOGIC_VECTOR(15 downto 0);
        y_421 : out STD_LOGIC_VECTOR(15 downto 0);
        y_422 : out STD_LOGIC_VECTOR(15 downto 0);
        y_423 : out STD_LOGIC_VECTOR(15 downto 0);
        y_424 : out STD_LOGIC_VECTOR(15 downto 0);
        y_425 : out STD_LOGIC_VECTOR(15 downto 0);
        y_426 : out STD_LOGIC_VECTOR(15 downto 0);
        y_427 : out STD_LOGIC_VECTOR(15 downto 0);
        y_428 : out STD_LOGIC_VECTOR(15 downto 0);
        y_429 : out STD_LOGIC_VECTOR(15 downto 0);
        y_430 : out STD_LOGIC_VECTOR(15 downto 0);
        y_431 : out STD_LOGIC_VECTOR(15 downto 0);
        y_432 : out STD_LOGIC_VECTOR(15 downto 0);
        y_433 : out STD_LOGIC_VECTOR(15 downto 0);
        y_434 : out STD_LOGIC_VECTOR(15 downto 0);
        y_435 : out STD_LOGIC_VECTOR(15 downto 0);
        y_436 : out STD_LOGIC_VECTOR(15 downto 0);
        y_437 : out STD_LOGIC_VECTOR(15 downto 0);
        y_438 : out STD_LOGIC_VECTOR(15 downto 0);
        y_439 : out STD_LOGIC_VECTOR(15 downto 0);
        y_440 : out STD_LOGIC_VECTOR(15 downto 0);
        y_441 : out STD_LOGIC_VECTOR(15 downto 0);
        y_442 : out STD_LOGIC_VECTOR(15 downto 0);
        y_443 : out STD_LOGIC_VECTOR(15 downto 0);
        y_444 : out STD_LOGIC_VECTOR(15 downto 0);
        y_445 : out STD_LOGIC_VECTOR(15 downto 0);
        y_446 : out STD_LOGIC_VECTOR(15 downto 0);
        y_447 : out STD_LOGIC_VECTOR(15 downto 0);
        y_448 : out STD_LOGIC_VECTOR(15 downto 0);
        y_449 : out STD_LOGIC_VECTOR(15 downto 0);
        y_450 : out STD_LOGIC_VECTOR(15 downto 0);
        y_451 : out STD_LOGIC_VECTOR(15 downto 0);
        y_452 : out STD_LOGIC_VECTOR(15 downto 0);
        y_453 : out STD_LOGIC_VECTOR(15 downto 0);
        y_454 : out STD_LOGIC_VECTOR(15 downto 0);
        y_455 : out STD_LOGIC_VECTOR(15 downto 0);
        y_456 : out STD_LOGIC_VECTOR(15 downto 0);
        y_457 : out STD_LOGIC_VECTOR(15 downto 0);
        y_458 : out STD_LOGIC_VECTOR(15 downto 0);
        y_459 : out STD_LOGIC_VECTOR(15 downto 0);
        y_460 : out STD_LOGIC_VECTOR(15 downto 0);
        y_461 : out STD_LOGIC_VECTOR(15 downto 0);
        y_462 : out STD_LOGIC_VECTOR(15 downto 0);
        y_463 : out STD_LOGIC_VECTOR(15 downto 0);
        y_464 : out STD_LOGIC_VECTOR(15 downto 0);
        y_465 : out STD_LOGIC_VECTOR(15 downto 0);
        y_466 : out STD_LOGIC_VECTOR(15 downto 0);
        y_467 : out STD_LOGIC_VECTOR(15 downto 0);
        y_468 : out STD_LOGIC_VECTOR(15 downto 0);
        y_469 : out STD_LOGIC_VECTOR(15 downto 0);
        y_470 : out STD_LOGIC_VECTOR(15 downto 0);
        y_471 : out STD_LOGIC_VECTOR(15 downto 0);
        y_472 : out STD_LOGIC_VECTOR(15 downto 0);
        y_473 : out STD_LOGIC_VECTOR(15 downto 0);
        y_474 : out STD_LOGIC_VECTOR(15 downto 0);
        y_475 : out STD_LOGIC_VECTOR(15 downto 0);
        y_476 : out STD_LOGIC_VECTOR(15 downto 0);
        y_477 : out STD_LOGIC_VECTOR(15 downto 0);
        y_478 : out STD_LOGIC_VECTOR(15 downto 0);
        y_479 : out STD_LOGIC_VECTOR(15 downto 0);
        y_480 : out STD_LOGIC_VECTOR(15 downto 0);
        y_481 : out STD_LOGIC_VECTOR(15 downto 0);
        y_482 : out STD_LOGIC_VECTOR(15 downto 0);
        y_483 : out STD_LOGIC_VECTOR(15 downto 0);
        y_484 : out STD_LOGIC_VECTOR(15 downto 0);
        y_485 : out STD_LOGIC_VECTOR(15 downto 0);
        y_486 : out STD_LOGIC_VECTOR(15 downto 0);
        y_487 : out STD_LOGIC_VECTOR(15 downto 0);
        y_488 : out STD_LOGIC_VECTOR(15 downto 0);
        y_489 : out STD_LOGIC_VECTOR(15 downto 0);
        y_490 : out STD_LOGIC_VECTOR(15 downto 0);
        y_491 : out STD_LOGIC_VECTOR(15 downto 0);
        y_492 : out STD_LOGIC_VECTOR(15 downto 0);
        y_493 : out STD_LOGIC_VECTOR(15 downto 0);
        y_494 : out STD_LOGIC_VECTOR(15 downto 0);
        y_495 : out STD_LOGIC_VECTOR(15 downto 0);
        y_496 : out STD_LOGIC_VECTOR(15 downto 0);
        y_497 : out STD_LOGIC_VECTOR(15 downto 0);
        y_498 : out STD_LOGIC_VECTOR(15 downto 0);
        y_499 : out STD_LOGIC_VECTOR(15 downto 0);
        y_500 : out STD_LOGIC_VECTOR(15 downto 0);
        y_501 : out STD_LOGIC_VECTOR(15 downto 0);
        y_502 : out STD_LOGIC_VECTOR(15 downto 0);
        y_503 : out STD_LOGIC_VECTOR(15 downto 0);
        y_504 : out STD_LOGIC_VECTOR(15 downto 0);
        y_505 : out STD_LOGIC_VECTOR(15 downto 0);
        y_506 : out STD_LOGIC_VECTOR(15 downto 0);
        y_507 : out STD_LOGIC_VECTOR(15 downto 0);
        y_508 : out STD_LOGIC_VECTOR(15 downto 0);
        y_509 : out STD_LOGIC_VECTOR(15 downto 0);
        y_510 : out STD_LOGIC_VECTOR(15 downto 0);
        y_511 : out STD_LOGIC_VECTOR(15 downto 0);
        y_512 : out STD_LOGIC_VECTOR(15 downto 0);
        y_513 : out STD_LOGIC_VECTOR(15 downto 0);
        y_514 : out STD_LOGIC_VECTOR(15 downto 0);
        y_515 : out STD_LOGIC_VECTOR(15 downto 0);
        y_516 : out STD_LOGIC_VECTOR(15 downto 0);
        y_517 : out STD_LOGIC_VECTOR(15 downto 0);
        y_518 : out STD_LOGIC_VECTOR(15 downto 0);
        y_519 : out STD_LOGIC_VECTOR(15 downto 0);
        y_520 : out STD_LOGIC_VECTOR(15 downto 0);
        y_521 : out STD_LOGIC_VECTOR(15 downto 0);
        y_522 : out STD_LOGIC_VECTOR(15 downto 0);
        y_523 : out STD_LOGIC_VECTOR(15 downto 0);
        y_524 : out STD_LOGIC_VECTOR(15 downto 0);
        y_525 : out STD_LOGIC_VECTOR(15 downto 0);
        y_526 : out STD_LOGIC_VECTOR(15 downto 0);
        y_527 : out STD_LOGIC_VECTOR(15 downto 0);
        y_528 : out STD_LOGIC_VECTOR(15 downto 0);
        y_529 : out STD_LOGIC_VECTOR(15 downto 0);
        y_530 : out STD_LOGIC_VECTOR(15 downto 0);
        y_531 : out STD_LOGIC_VECTOR(15 downto 0);
        y_532 : out STD_LOGIC_VECTOR(15 downto 0);
        y_533 : out STD_LOGIC_VECTOR(15 downto 0);
        y_534 : out STD_LOGIC_VECTOR(15 downto 0);
        y_535 : out STD_LOGIC_VECTOR(15 downto 0);
        y_536 : out STD_LOGIC_VECTOR(15 downto 0);
        y_537 : out STD_LOGIC_VECTOR(15 downto 0);
        y_538 : out STD_LOGIC_VECTOR(15 downto 0);
        y_539 : out STD_LOGIC_VECTOR(15 downto 0);
        y_540 : out STD_LOGIC_VECTOR(15 downto 0);
        y_541 : out STD_LOGIC_VECTOR(15 downto 0);
        y_542 : out STD_LOGIC_VECTOR(15 downto 0);
        y_543 : out STD_LOGIC_VECTOR(15 downto 0);
        y_544 : out STD_LOGIC_VECTOR(15 downto 0);
        y_545 : out STD_LOGIC_VECTOR(15 downto 0);
        y_546 : out STD_LOGIC_VECTOR(15 downto 0);
        y_547 : out STD_LOGIC_VECTOR(15 downto 0);
        y_548 : out STD_LOGIC_VECTOR(15 downto 0);
        y_549 : out STD_LOGIC_VECTOR(15 downto 0);
        y_550 : out STD_LOGIC_VECTOR(15 downto 0);
        y_551 : out STD_LOGIC_VECTOR(15 downto 0);
        y_552 : out STD_LOGIC_VECTOR(15 downto 0);
        y_553 : out STD_LOGIC_VECTOR(15 downto 0);
        y_554 : out STD_LOGIC_VECTOR(15 downto 0);
        y_555 : out STD_LOGIC_VECTOR(15 downto 0);
        y_556 : out STD_LOGIC_VECTOR(15 downto 0);
        y_557 : out STD_LOGIC_VECTOR(15 downto 0);
        y_558 : out STD_LOGIC_VECTOR(15 downto 0);
        y_559 : out STD_LOGIC_VECTOR(15 downto 0);
        y_560 : out STD_LOGIC_VECTOR(15 downto 0);
        y_561 : out STD_LOGIC_VECTOR(15 downto 0);
        y_562 : out STD_LOGIC_VECTOR(15 downto 0);
        y_563 : out STD_LOGIC_VECTOR(15 downto 0);
        y_564 : out STD_LOGIC_VECTOR(15 downto 0);
        y_565 : out STD_LOGIC_VECTOR(15 downto 0);
        y_566 : out STD_LOGIC_VECTOR(15 downto 0);
        y_567 : out STD_LOGIC_VECTOR(15 downto 0);
        y_568 : out STD_LOGIC_VECTOR(15 downto 0);
        y_569 : out STD_LOGIC_VECTOR(15 downto 0);
        y_570 : out STD_LOGIC_VECTOR(15 downto 0);
        y_571 : out STD_LOGIC_VECTOR(15 downto 0);
        y_572 : out STD_LOGIC_VECTOR(15 downto 0);
        y_573 : out STD_LOGIC_VECTOR(15 downto 0);
        y_574 : out STD_LOGIC_VECTOR(15 downto 0);
        y_575 : out STD_LOGIC_VECTOR(15 downto 0);
        y_576 : out STD_LOGIC_VECTOR(15 downto 0);
        y_577 : out STD_LOGIC_VECTOR(15 downto 0);
        y_578 : out STD_LOGIC_VECTOR(15 downto 0);
        y_579 : out STD_LOGIC_VECTOR(15 downto 0);
        y_580 : out STD_LOGIC_VECTOR(15 downto 0);
        y_581 : out STD_LOGIC_VECTOR(15 downto 0);
        y_582 : out STD_LOGIC_VECTOR(15 downto 0);
        y_583 : out STD_LOGIC_VECTOR(15 downto 0);
        y_584 : out STD_LOGIC_VECTOR(15 downto 0);
        y_585 : out STD_LOGIC_VECTOR(15 downto 0);
        y_586 : out STD_LOGIC_VECTOR(15 downto 0);
        y_587 : out STD_LOGIC_VECTOR(15 downto 0);
        y_588 : out STD_LOGIC_VECTOR(15 downto 0);
        y_589 : out STD_LOGIC_VECTOR(15 downto 0);
        y_590 : out STD_LOGIC_VECTOR(15 downto 0);
        y_591 : out STD_LOGIC_VECTOR(15 downto 0);
        y_592 : out STD_LOGIC_VECTOR(15 downto 0);
        y_593 : out STD_LOGIC_VECTOR(15 downto 0);
        y_594 : out STD_LOGIC_VECTOR(15 downto 0);
        y_595 : out STD_LOGIC_VECTOR(15 downto 0);
        y_596 : out STD_LOGIC_VECTOR(15 downto 0);
        y_597 : out STD_LOGIC_VECTOR(15 downto 0);
        y_598 : out STD_LOGIC_VECTOR(15 downto 0);
        y_599 : out STD_LOGIC_VECTOR(15 downto 0);
        y_600 : out STD_LOGIC_VECTOR(15 downto 0);
        y_601 : out STD_LOGIC_VECTOR(15 downto 0);
        y_602 : out STD_LOGIC_VECTOR(15 downto 0);
        y_603 : out STD_LOGIC_VECTOR(15 downto 0);
        y_604 : out STD_LOGIC_VECTOR(15 downto 0);
        y_605 : out STD_LOGIC_VECTOR(15 downto 0);
        y_606 : out STD_LOGIC_VECTOR(15 downto 0);
        y_607 : out STD_LOGIC_VECTOR(15 downto 0);
        y_608 : out STD_LOGIC_VECTOR(15 downto 0);
        y_609 : out STD_LOGIC_VECTOR(15 downto 0);
        y_610 : out STD_LOGIC_VECTOR(15 downto 0);
        y_611 : out STD_LOGIC_VECTOR(15 downto 0);
        y_612 : out STD_LOGIC_VECTOR(15 downto 0);
        y_613 : out STD_LOGIC_VECTOR(15 downto 0);
        y_614 : out STD_LOGIC_VECTOR(15 downto 0);
        y_615 : out STD_LOGIC_VECTOR(15 downto 0);
        y_616 : out STD_LOGIC_VECTOR(15 downto 0);
        y_617 : out STD_LOGIC_VECTOR(15 downto 0);
        y_618 : out STD_LOGIC_VECTOR(15 downto 0);
        y_619 : out STD_LOGIC_VECTOR(15 downto 0);
        y_620 : out STD_LOGIC_VECTOR(15 downto 0);
        y_621 : out STD_LOGIC_VECTOR(15 downto 0);
        y_622 : out STD_LOGIC_VECTOR(15 downto 0);
        y_623 : out STD_LOGIC_VECTOR(15 downto 0);
        y_624 : out STD_LOGIC_VECTOR(15 downto 0);
        y_625 : out STD_LOGIC_VECTOR(15 downto 0);
        y_626 : out STD_LOGIC_VECTOR(15 downto 0);
        y_627 : out STD_LOGIC_VECTOR(15 downto 0);
        y_628 : out STD_LOGIC_VECTOR(15 downto 0);
        y_629 : out STD_LOGIC_VECTOR(15 downto 0);
        y_630 : out STD_LOGIC_VECTOR(15 downto 0);
        y_631 : out STD_LOGIC_VECTOR(15 downto 0);
        y_632 : out STD_LOGIC_VECTOR(15 downto 0);
        y_633 : out STD_LOGIC_VECTOR(15 downto 0);
        y_634 : out STD_LOGIC_VECTOR(15 downto 0);
        y_635 : out STD_LOGIC_VECTOR(15 downto 0);
        y_636 : out STD_LOGIC_VECTOR(15 downto 0);
        y_637 : out STD_LOGIC_VECTOR(15 downto 0);
        y_638 : out STD_LOGIC_VECTOR(15 downto 0);
        y_639 : out STD_LOGIC_VECTOR(15 downto 0);
        y_640 : out STD_LOGIC_VECTOR(15 downto 0);
        y_641 : out STD_LOGIC_VECTOR(15 downto 0);
        y_642 : out STD_LOGIC_VECTOR(15 downto 0);
        y_643 : out STD_LOGIC_VECTOR(15 downto 0);
        y_644 : out STD_LOGIC_VECTOR(15 downto 0);
        y_645 : out STD_LOGIC_VECTOR(15 downto 0);
        y_646 : out STD_LOGIC_VECTOR(15 downto 0);
        y_647 : out STD_LOGIC_VECTOR(15 downto 0);
        y_648 : out STD_LOGIC_VECTOR(15 downto 0);
        y_649 : out STD_LOGIC_VECTOR(15 downto 0);
        y_650 : out STD_LOGIC_VECTOR(15 downto 0);
        y_651 : out STD_LOGIC_VECTOR(15 downto 0);
        y_652 : out STD_LOGIC_VECTOR(15 downto 0);
        y_653 : out STD_LOGIC_VECTOR(15 downto 0);
        y_654 : out STD_LOGIC_VECTOR(15 downto 0);
        y_655 : out STD_LOGIC_VECTOR(15 downto 0);
        y_656 : out STD_LOGIC_VECTOR(15 downto 0);
        y_657 : out STD_LOGIC_VECTOR(15 downto 0);
        y_658 : out STD_LOGIC_VECTOR(15 downto 0);
        y_659 : out STD_LOGIC_VECTOR(15 downto 0);
        y_660 : out STD_LOGIC_VECTOR(15 downto 0);
        y_661 : out STD_LOGIC_VECTOR(15 downto 0);
        y_662 : out STD_LOGIC_VECTOR(15 downto 0);
        y_663 : out STD_LOGIC_VECTOR(15 downto 0);
        y_664 : out STD_LOGIC_VECTOR(15 downto 0);
        y_665 : out STD_LOGIC_VECTOR(15 downto 0);
        y_666 : out STD_LOGIC_VECTOR(15 downto 0);
        y_667 : out STD_LOGIC_VECTOR(15 downto 0);
        y_668 : out STD_LOGIC_VECTOR(15 downto 0);
        y_669 : out STD_LOGIC_VECTOR(15 downto 0);
        y_670 : out STD_LOGIC_VECTOR(15 downto 0);
        y_671 : out STD_LOGIC_VECTOR(15 downto 0);
        y_672 : out STD_LOGIC_VECTOR(15 downto 0);
        y_673 : out STD_LOGIC_VECTOR(15 downto 0);
        y_674 : out STD_LOGIC_VECTOR(15 downto 0);
        y_675 : out STD_LOGIC_VECTOR(15 downto 0);
        y_676 : out STD_LOGIC_VECTOR(15 downto 0);
        y_677 : out STD_LOGIC_VECTOR(15 downto 0);
        y_678 : out STD_LOGIC_VECTOR(15 downto 0);
        y_679 : out STD_LOGIC_VECTOR(15 downto 0);
        y_680 : out STD_LOGIC_VECTOR(15 downto 0);
        y_681 : out STD_LOGIC_VECTOR(15 downto 0);
        y_682 : out STD_LOGIC_VECTOR(15 downto 0);
        y_683 : out STD_LOGIC_VECTOR(15 downto 0);
        y_684 : out STD_LOGIC_VECTOR(15 downto 0);
        y_685 : out STD_LOGIC_VECTOR(15 downto 0);
        y_686 : out STD_LOGIC_VECTOR(15 downto 0);
        y_687 : out STD_LOGIC_VECTOR(15 downto 0);
        y_688 : out STD_LOGIC_VECTOR(15 downto 0);
        y_689 : out STD_LOGIC_VECTOR(15 downto 0);
        y_690 : out STD_LOGIC_VECTOR(15 downto 0);
        y_691 : out STD_LOGIC_VECTOR(15 downto 0);
        y_692 : out STD_LOGIC_VECTOR(15 downto 0);
        y_693 : out STD_LOGIC_VECTOR(15 downto 0);
        y_694 : out STD_LOGIC_VECTOR(15 downto 0);
        y_695 : out STD_LOGIC_VECTOR(15 downto 0);
        y_696 : out STD_LOGIC_VECTOR(15 downto 0);
        y_697 : out STD_LOGIC_VECTOR(15 downto 0);
        y_698 : out STD_LOGIC_VECTOR(15 downto 0);
        y_699 : out STD_LOGIC_VECTOR(15 downto 0);
        y_700 : out STD_LOGIC_VECTOR(15 downto 0);
        y_701 : out STD_LOGIC_VECTOR(15 downto 0);
        y_702 : out STD_LOGIC_VECTOR(15 downto 0);
        y_703 : out STD_LOGIC_VECTOR(15 downto 0);
        y_704 : out STD_LOGIC_VECTOR(15 downto 0);
        y_705 : out STD_LOGIC_VECTOR(15 downto 0);
        y_706 : out STD_LOGIC_VECTOR(15 downto 0);
        y_707 : out STD_LOGIC_VECTOR(15 downto 0);
        y_708 : out STD_LOGIC_VECTOR(15 downto 0);
        y_709 : out STD_LOGIC_VECTOR(15 downto 0);
        y_710 : out STD_LOGIC_VECTOR(15 downto 0);
        y_711 : out STD_LOGIC_VECTOR(15 downto 0);
        y_712 : out STD_LOGIC_VECTOR(15 downto 0);
        y_713 : out STD_LOGIC_VECTOR(15 downto 0);
        y_714 : out STD_LOGIC_VECTOR(15 downto 0);
        y_715 : out STD_LOGIC_VECTOR(15 downto 0);
        y_716 : out STD_LOGIC_VECTOR(15 downto 0);
        y_717 : out STD_LOGIC_VECTOR(15 downto 0);
        y_718 : out STD_LOGIC_VECTOR(15 downto 0);
        y_719 : out STD_LOGIC_VECTOR(15 downto 0);
        y_720 : out STD_LOGIC_VECTOR(15 downto 0);
        y_721 : out STD_LOGIC_VECTOR(15 downto 0);
        y_722 : out STD_LOGIC_VECTOR(15 downto 0);
        y_723 : out STD_LOGIC_VECTOR(15 downto 0);
        y_724 : out STD_LOGIC_VECTOR(15 downto 0);
        y_725 : out STD_LOGIC_VECTOR(15 downto 0);
        y_726 : out STD_LOGIC_VECTOR(15 downto 0);
        y_727 : out STD_LOGIC_VECTOR(15 downto 0);
        y_728 : out STD_LOGIC_VECTOR(15 downto 0);
        y_729 : out STD_LOGIC_VECTOR(15 downto 0);
        y_730 : out STD_LOGIC_VECTOR(15 downto 0);
        y_731 : out STD_LOGIC_VECTOR(15 downto 0);
        y_732 : out STD_LOGIC_VECTOR(15 downto 0);
        y_733 : out STD_LOGIC_VECTOR(15 downto 0);
        y_734 : out STD_LOGIC_VECTOR(15 downto 0);
        y_735 : out STD_LOGIC_VECTOR(15 downto 0);
        y_736 : out STD_LOGIC_VECTOR(15 downto 0);
        y_737 : out STD_LOGIC_VECTOR(15 downto 0);
        y_738 : out STD_LOGIC_VECTOR(15 downto 0);
        y_739 : out STD_LOGIC_VECTOR(15 downto 0);
        y_740 : out STD_LOGIC_VECTOR(15 downto 0);
        y_741 : out STD_LOGIC_VECTOR(15 downto 0);
        y_742 : out STD_LOGIC_VECTOR(15 downto 0);
        y_743 : out STD_LOGIC_VECTOR(15 downto 0);
        y_744 : out STD_LOGIC_VECTOR(15 downto 0);
        y_745 : out STD_LOGIC_VECTOR(15 downto 0);
        y_746 : out STD_LOGIC_VECTOR(15 downto 0);
        y_747 : out STD_LOGIC_VECTOR(15 downto 0);
        y_748 : out STD_LOGIC_VECTOR(15 downto 0);
        y_749 : out STD_LOGIC_VECTOR(15 downto 0);
        y_750 : out STD_LOGIC_VECTOR(15 downto 0);
        y_751 : out STD_LOGIC_VECTOR(15 downto 0);
        y_752 : out STD_LOGIC_VECTOR(15 downto 0);
        y_753 : out STD_LOGIC_VECTOR(15 downto 0);
        y_754 : out STD_LOGIC_VECTOR(15 downto 0);
        y_755 : out STD_LOGIC_VECTOR(15 downto 0);
        y_756 : out STD_LOGIC_VECTOR(15 downto 0);
        y_757 : out STD_LOGIC_VECTOR(15 downto 0);
        y_758 : out STD_LOGIC_VECTOR(15 downto 0);
        y_759 : out STD_LOGIC_VECTOR(15 downto 0);
        y_760 : out STD_LOGIC_VECTOR(15 downto 0);
        y_761 : out STD_LOGIC_VECTOR(15 downto 0);
        y_762 : out STD_LOGIC_VECTOR(15 downto 0);
        y_763 : out STD_LOGIC_VECTOR(15 downto 0);
        y_764 : out STD_LOGIC_VECTOR(15 downto 0);
        y_765 : out STD_LOGIC_VECTOR(15 downto 0);
        y_766 : out STD_LOGIC_VECTOR(15 downto 0);
        y_767 : out STD_LOGIC_VECTOR(15 downto 0);
        y_768 : out STD_LOGIC_VECTOR(15 downto 0);
        y_769 : out STD_LOGIC_VECTOR(15 downto 0);
        y_770 : out STD_LOGIC_VECTOR(15 downto 0);
        y_771 : out STD_LOGIC_VECTOR(15 downto 0);
        y_772 : out STD_LOGIC_VECTOR(15 downto 0);
        y_773 : out STD_LOGIC_VECTOR(15 downto 0);
        y_774 : out STD_LOGIC_VECTOR(15 downto 0);
        y_775 : out STD_LOGIC_VECTOR(15 downto 0);
        y_776 : out STD_LOGIC_VECTOR(15 downto 0);
        y_777 : out STD_LOGIC_VECTOR(15 downto 0);
        y_778 : out STD_LOGIC_VECTOR(15 downto 0);
        y_779 : out STD_LOGIC_VECTOR(15 downto 0);
        y_780 : out STD_LOGIC_VECTOR(15 downto 0);
        y_781 : out STD_LOGIC_VECTOR(15 downto 0);
        y_782 : out STD_LOGIC_VECTOR(15 downto 0);
        y_783 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end lstm_layer ;
architecture Behavioral of lstm_layer is

component lstm_layer_4 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_4;
component lstm_layer_5 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_5;
component lstm_layer_6 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_6;
component lstm_layer_7 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_7;
component lstm_layer_8 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_8;
component lstm_layer_9 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_9;
component lstm_layer_10 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_10;
component lstm_layer_11 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_11;
component lstm_layer_12 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_12;
component lstm_layer_13 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_13;
component lstm_layer_14 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_14;
component lstm_layer_15 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_15;
component lstm_layer_16 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_16;
component lstm_layer_17 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_17;
component lstm_layer_18 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_18;
component lstm_layer_19 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_19;
component lstm_layer_20 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_20;
component lstm_layer_21 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_21;
component lstm_layer_22 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_22;
component lstm_layer_23 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_23;
component lstm_layer_24 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_24;
component lstm_layer_25 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_25;
component lstm_layer_26 is
	Port (
		 x_0 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_1 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_2 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_3 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_4 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_5 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_6 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_7 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_8 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_9 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_10 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_11 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_12 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_13 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_14 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_15 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_16 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_17 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_18 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_19 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_20 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_21 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_22 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_23 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_24 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_25 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_26 : in STD_LOGIC_VECTOR(15 downto 0);
		 x_27 : in STD_LOGIC_VECTOR(15 downto 0);
		 y_0 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_1 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_2 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_3 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_4 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_5 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_6 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_7 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_8 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_9 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_10 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_11 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_12 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_13 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_14 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_15 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_16 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_17 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_18 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_19 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_20 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_21 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_22 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_23 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_24 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_25 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_26 : out STD_LOGIC_VECTOR(15 downto 0);
		 y_27 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component lstm_layer_26;

begin

ut4_lstm_layer_4: lstm_layer_4 port map(
	x_0 => x_112,
	x_1 => x_113,
	x_2 => x_114,
	x_3 => x_115,
	x_4 => x_116,
	x_5 => x_117,
	x_6 => x_118,
	x_7 => x_119,
	x_8 => x_120,
	x_9 => x_121,
	x_10 => x_122,
	x_11 => x_123,
	x_12 => x_124,
	x_13 => x_125,
	x_14 => x_126,
	x_15 => x_127,
	x_16 => x_128,
	x_17 => x_129,
	x_18 => x_130,
	x_19 => x_131,
	x_20 => x_132,
	x_21 => x_133,
	x_22 => x_134,
	x_23 => x_135,
	x_24 => x_136,
	x_25 => x_137,
	x_26 => x_138,
	x_27 => x_139,
	y_0 => y_112,
	y_1 => y_113,
	y_2 => y_114,
	y_3 => y_115,
	y_4 => y_116,
	y_5 => y_117,
	y_6 => y_118,
	y_7 => y_119,
	y_8 => y_120,
	y_9 => y_121,
	y_10 => y_122,
	y_11 => y_123,
	y_12 => y_124,
	y_13 => y_125,
	y_14 => y_126,
	y_15 => y_127,
	y_16 => y_128,
	y_17 => y_129,
	y_18 => y_130,
	y_19 => y_131,
	y_20 => y_132,
	y_21 => y_133,
	y_22 => y_134,
	y_23 => y_135,
	y_24 => y_136,
	y_25 => y_137,
	y_26 => y_138,
	y_27 => y_139
    );
ut5_lstm_layer_5: lstm_layer_5 port map(
	x_0 => x_140,
	x_1 => x_141,
	x_2 => x_142,
	x_3 => x_143,
	x_4 => x_144,
	x_5 => x_145,
	x_6 => x_146,
	x_7 => x_147,
	x_8 => x_148,
	x_9 => x_149,
	x_10 => x_150,
	x_11 => x_151,
	x_12 => x_152,
	x_13 => x_153,
	x_14 => x_154,
	x_15 => x_155,
	x_16 => x_156,
	x_17 => x_157,
	x_18 => x_158,
	x_19 => x_159,
	x_20 => x_160,
	x_21 => x_161,
	x_22 => x_162,
	x_23 => x_163,
	x_24 => x_164,
	x_25 => x_165,
	x_26 => x_166,
	x_27 => x_167,
	y_0 => y_140,
	y_1 => y_141,
	y_2 => y_142,
	y_3 => y_143,
	y_4 => y_144,
	y_5 => y_145,
	y_6 => y_146,
	y_7 => y_147,
	y_8 => y_148,
	y_9 => y_149,
	y_10 => y_150,
	y_11 => y_151,
	y_12 => y_152,
	y_13 => y_153,
	y_14 => y_154,
	y_15 => y_155,
	y_16 => y_156,
	y_17 => y_157,
	y_18 => y_158,
	y_19 => y_159,
	y_20 => y_160,
	y_21 => y_161,
	y_22 => y_162,
	y_23 => y_163,
	y_24 => y_164,
	y_25 => y_165,
	y_26 => y_166,
	y_27 => y_167
    );
ut6_lstm_layer_6: lstm_layer_6 port map(
	x_0 => x_168,
	x_1 => x_169,
	x_2 => x_170,
	x_3 => x_171,
	x_4 => x_172,
	x_5 => x_173,
	x_6 => x_174,
	x_7 => x_175,
	x_8 => x_176,
	x_9 => x_177,
	x_10 => x_178,
	x_11 => x_179,
	x_12 => x_180,
	x_13 => x_181,
	x_14 => x_182,
	x_15 => x_183,
	x_16 => x_184,
	x_17 => x_185,
	x_18 => x_186,
	x_19 => x_187,
	x_20 => x_188,
	x_21 => x_189,
	x_22 => x_190,
	x_23 => x_191,
	x_24 => x_192,
	x_25 => x_193,
	x_26 => x_194,
	x_27 => x_195,
	y_0 => y_168,
	y_1 => y_169,
	y_2 => y_170,
	y_3 => y_171,
	y_4 => y_172,
	y_5 => y_173,
	y_6 => y_174,
	y_7 => y_175,
	y_8 => y_176,
	y_9 => y_177,
	y_10 => y_178,
	y_11 => y_179,
	y_12 => y_180,
	y_13 => y_181,
	y_14 => y_182,
	y_15 => y_183,
	y_16 => y_184,
	y_17 => y_185,
	y_18 => y_186,
	y_19 => y_187,
	y_20 => y_188,
	y_21 => y_189,
	y_22 => y_190,
	y_23 => y_191,
	y_24 => y_192,
	y_25 => y_193,
	y_26 => y_194,
	y_27 => y_195
    );
ut7_lstm_layer_7: lstm_layer_7 port map(
	x_0 => x_196,
	x_1 => x_197,
	x_2 => x_198,
	x_3 => x_199,
	x_4 => x_200,
	x_5 => x_201,
	x_6 => x_202,
	x_7 => x_203,
	x_8 => x_204,
	x_9 => x_205,
	x_10 => x_206,
	x_11 => x_207,
	x_12 => x_208,
	x_13 => x_209,
	x_14 => x_210,
	x_15 => x_211,
	x_16 => x_212,
	x_17 => x_213,
	x_18 => x_214,
	x_19 => x_215,
	x_20 => x_216,
	x_21 => x_217,
	x_22 => x_218,
	x_23 => x_219,
	x_24 => x_220,
	x_25 => x_221,
	x_26 => x_222,
	x_27 => x_223,
	y_0 => y_196,
	y_1 => y_197,
	y_2 => y_198,
	y_3 => y_199,
	y_4 => y_200,
	y_5 => y_201,
	y_6 => y_202,
	y_7 => y_203,
	y_8 => y_204,
	y_9 => y_205,
	y_10 => y_206,
	y_11 => y_207,
	y_12 => y_208,
	y_13 => y_209,
	y_14 => y_210,
	y_15 => y_211,
	y_16 => y_212,
	y_17 => y_213,
	y_18 => y_214,
	y_19 => y_215,
	y_20 => y_216,
	y_21 => y_217,
	y_22 => y_218,
	y_23 => y_219,
	y_24 => y_220,
	y_25 => y_221,
	y_26 => y_222,
	y_27 => y_223
    );
ut8_lstm_layer_8: lstm_layer_8 port map(
	x_0 => x_224,
	x_1 => x_225,
	x_2 => x_226,
	x_3 => x_227,
	x_4 => x_228,
	x_5 => x_229,
	x_6 => x_230,
	x_7 => x_231,
	x_8 => x_232,
	x_9 => x_233,
	x_10 => x_234,
	x_11 => x_235,
	x_12 => x_236,
	x_13 => x_237,
	x_14 => x_238,
	x_15 => x_239,
	x_16 => x_240,
	x_17 => x_241,
	x_18 => x_242,
	x_19 => x_243,
	x_20 => x_244,
	x_21 => x_245,
	x_22 => x_246,
	x_23 => x_247,
	x_24 => x_248,
	x_25 => x_249,
	x_26 => x_250,
	x_27 => x_251,
	y_0 => y_224,
	y_1 => y_225,
	y_2 => y_226,
	y_3 => y_227,
	y_4 => y_228,
	y_5 => y_229,
	y_6 => y_230,
	y_7 => y_231,
	y_8 => y_232,
	y_9 => y_233,
	y_10 => y_234,
	y_11 => y_235,
	y_12 => y_236,
	y_13 => y_237,
	y_14 => y_238,
	y_15 => y_239,
	y_16 => y_240,
	y_17 => y_241,
	y_18 => y_242,
	y_19 => y_243,
	y_20 => y_244,
	y_21 => y_245,
	y_22 => y_246,
	y_23 => y_247,
	y_24 => y_248,
	y_25 => y_249,
	y_26 => y_250,
	y_27 => y_251
    );
ut9_lstm_layer_9: lstm_layer_9 port map(
	x_0 => x_252,
	x_1 => x_253,
	x_2 => x_254,
	x_3 => x_255,
	x_4 => x_256,
	x_5 => x_257,
	x_6 => x_258,
	x_7 => x_259,
	x_8 => x_260,
	x_9 => x_261,
	x_10 => x_262,
	x_11 => x_263,
	x_12 => x_264,
	x_13 => x_265,
	x_14 => x_266,
	x_15 => x_267,
	x_16 => x_268,
	x_17 => x_269,
	x_18 => x_270,
	x_19 => x_271,
	x_20 => x_272,
	x_21 => x_273,
	x_22 => x_274,
	x_23 => x_275,
	x_24 => x_276,
	x_25 => x_277,
	x_26 => x_278,
	x_27 => x_279,
	y_0 => y_252,
	y_1 => y_253,
	y_2 => y_254,
	y_3 => y_255,
	y_4 => y_256,
	y_5 => y_257,
	y_6 => y_258,
	y_7 => y_259,
	y_8 => y_260,
	y_9 => y_261,
	y_10 => y_262,
	y_11 => y_263,
	y_12 => y_264,
	y_13 => y_265,
	y_14 => y_266,
	y_15 => y_267,
	y_16 => y_268,
	y_17 => y_269,
	y_18 => y_270,
	y_19 => y_271,
	y_20 => y_272,
	y_21 => y_273,
	y_22 => y_274,
	y_23 => y_275,
	y_24 => y_276,
	y_25 => y_277,
	y_26 => y_278,
	y_27 => y_279
    );
ut10_lstm_layer_10: lstm_layer_10 port map(
	x_0 => x_280,
	x_1 => x_281,
	x_2 => x_282,
	x_3 => x_283,
	x_4 => x_284,
	x_5 => x_285,
	x_6 => x_286,
	x_7 => x_287,
	x_8 => x_288,
	x_9 => x_289,
	x_10 => x_290,
	x_11 => x_291,
	x_12 => x_292,
	x_13 => x_293,
	x_14 => x_294,
	x_15 => x_295,
	x_16 => x_296,
	x_17 => x_297,
	x_18 => x_298,
	x_19 => x_299,
	x_20 => x_300,
	x_21 => x_301,
	x_22 => x_302,
	x_23 => x_303,
	x_24 => x_304,
	x_25 => x_305,
	x_26 => x_306,
	x_27 => x_307,
	y_0 => y_280,
	y_1 => y_281,
	y_2 => y_282,
	y_3 => y_283,
	y_4 => y_284,
	y_5 => y_285,
	y_6 => y_286,
	y_7 => y_287,
	y_8 => y_288,
	y_9 => y_289,
	y_10 => y_290,
	y_11 => y_291,
	y_12 => y_292,
	y_13 => y_293,
	y_14 => y_294,
	y_15 => y_295,
	y_16 => y_296,
	y_17 => y_297,
	y_18 => y_298,
	y_19 => y_299,
	y_20 => y_300,
	y_21 => y_301,
	y_22 => y_302,
	y_23 => y_303,
	y_24 => y_304,
	y_25 => y_305,
	y_26 => y_306,
	y_27 => y_307
    );
ut11_lstm_layer_11: lstm_layer_11 port map(
	x_0 => x_308,
	x_1 => x_309,
	x_2 => x_310,
	x_3 => x_311,
	x_4 => x_312,
	x_5 => x_313,
	x_6 => x_314,
	x_7 => x_315,
	x_8 => x_316,
	x_9 => x_317,
	x_10 => x_318,
	x_11 => x_319,
	x_12 => x_320,
	x_13 => x_321,
	x_14 => x_322,
	x_15 => x_323,
	x_16 => x_324,
	x_17 => x_325,
	x_18 => x_326,
	x_19 => x_327,
	x_20 => x_328,
	x_21 => x_329,
	x_22 => x_330,
	x_23 => x_331,
	x_24 => x_332,
	x_25 => x_333,
	x_26 => x_334,
	x_27 => x_335,
	y_0 => y_308,
	y_1 => y_309,
	y_2 => y_310,
	y_3 => y_311,
	y_4 => y_312,
	y_5 => y_313,
	y_6 => y_314,
	y_7 => y_315,
	y_8 => y_316,
	y_9 => y_317,
	y_10 => y_318,
	y_11 => y_319,
	y_12 => y_320,
	y_13 => y_321,
	y_14 => y_322,
	y_15 => y_323,
	y_16 => y_324,
	y_17 => y_325,
	y_18 => y_326,
	y_19 => y_327,
	y_20 => y_328,
	y_21 => y_329,
	y_22 => y_330,
	y_23 => y_331,
	y_24 => y_332,
	y_25 => y_333,
	y_26 => y_334,
	y_27 => y_335
    );
ut12_lstm_layer_12: lstm_layer_12 port map(
	x_0 => x_336,
	x_1 => x_337,
	x_2 => x_338,
	x_3 => x_339,
	x_4 => x_340,
	x_5 => x_341,
	x_6 => x_342,
	x_7 => x_343,
	x_8 => x_344,
	x_9 => x_345,
	x_10 => x_346,
	x_11 => x_347,
	x_12 => x_348,
	x_13 => x_349,
	x_14 => x_350,
	x_15 => x_351,
	x_16 => x_352,
	x_17 => x_353,
	x_18 => x_354,
	x_19 => x_355,
	x_20 => x_356,
	x_21 => x_357,
	x_22 => x_358,
	x_23 => x_359,
	x_24 => x_360,
	x_25 => x_361,
	x_26 => x_362,
	x_27 => x_363,
	y_0 => y_336,
	y_1 => y_337,
	y_2 => y_338,
	y_3 => y_339,
	y_4 => y_340,
	y_5 => y_341,
	y_6 => y_342,
	y_7 => y_343,
	y_8 => y_344,
	y_9 => y_345,
	y_10 => y_346,
	y_11 => y_347,
	y_12 => y_348,
	y_13 => y_349,
	y_14 => y_350,
	y_15 => y_351,
	y_16 => y_352,
	y_17 => y_353,
	y_18 => y_354,
	y_19 => y_355,
	y_20 => y_356,
	y_21 => y_357,
	y_22 => y_358,
	y_23 => y_359,
	y_24 => y_360,
	y_25 => y_361,
	y_26 => y_362,
	y_27 => y_363
    );
ut13_lstm_layer_13: lstm_layer_13 port map(
	x_0 => x_364,
	x_1 => x_365,
	x_2 => x_366,
	x_3 => x_367,
	x_4 => x_368,
	x_5 => x_369,
	x_6 => x_370,
	x_7 => x_371,
	x_8 => x_372,
	x_9 => x_373,
	x_10 => x_374,
	x_11 => x_375,
	x_12 => x_376,
	x_13 => x_377,
	x_14 => x_378,
	x_15 => x_379,
	x_16 => x_380,
	x_17 => x_381,
	x_18 => x_382,
	x_19 => x_383,
	x_20 => x_384,
	x_21 => x_385,
	x_22 => x_386,
	x_23 => x_387,
	x_24 => x_388,
	x_25 => x_389,
	x_26 => x_390,
	x_27 => x_391,
	y_0 => y_364,
	y_1 => y_365,
	y_2 => y_366,
	y_3 => y_367,
	y_4 => y_368,
	y_5 => y_369,
	y_6 => y_370,
	y_7 => y_371,
	y_8 => y_372,
	y_9 => y_373,
	y_10 => y_374,
	y_11 => y_375,
	y_12 => y_376,
	y_13 => y_377,
	y_14 => y_378,
	y_15 => y_379,
	y_16 => y_380,
	y_17 => y_381,
	y_18 => y_382,
	y_19 => y_383,
	y_20 => y_384,
	y_21 => y_385,
	y_22 => y_386,
	y_23 => y_387,
	y_24 => y_388,
	y_25 => y_389,
	y_26 => y_390,
	y_27 => y_391
    );
ut14_lstm_layer_14: lstm_layer_14 port map(
	x_0 => x_392,
	x_1 => x_393,
	x_2 => x_394,
	x_3 => x_395,
	x_4 => x_396,
	x_5 => x_397,
	x_6 => x_398,
	x_7 => x_399,
	x_8 => x_400,
	x_9 => x_401,
	x_10 => x_402,
	x_11 => x_403,
	x_12 => x_404,
	x_13 => x_405,
	x_14 => x_406,
	x_15 => x_407,
	x_16 => x_408,
	x_17 => x_409,
	x_18 => x_410,
	x_19 => x_411,
	x_20 => x_412,
	x_21 => x_413,
	x_22 => x_414,
	x_23 => x_415,
	x_24 => x_416,
	x_25 => x_417,
	x_26 => x_418,
	x_27 => x_419,
	y_0 => y_392,
	y_1 => y_393,
	y_2 => y_394,
	y_3 => y_395,
	y_4 => y_396,
	y_5 => y_397,
	y_6 => y_398,
	y_7 => y_399,
	y_8 => y_400,
	y_9 => y_401,
	y_10 => y_402,
	y_11 => y_403,
	y_12 => y_404,
	y_13 => y_405,
	y_14 => y_406,
	y_15 => y_407,
	y_16 => y_408,
	y_17 => y_409,
	y_18 => y_410,
	y_19 => y_411,
	y_20 => y_412,
	y_21 => y_413,
	y_22 => y_414,
	y_23 => y_415,
	y_24 => y_416,
	y_25 => y_417,
	y_26 => y_418,
	y_27 => y_419
    );
ut15_lstm_layer_15: lstm_layer_15 port map(
	x_0 => x_420,
	x_1 => x_421,
	x_2 => x_422,
	x_3 => x_423,
	x_4 => x_424,
	x_5 => x_425,
	x_6 => x_426,
	x_7 => x_427,
	x_8 => x_428,
	x_9 => x_429,
	x_10 => x_430,
	x_11 => x_431,
	x_12 => x_432,
	x_13 => x_433,
	x_14 => x_434,
	x_15 => x_435,
	x_16 => x_436,
	x_17 => x_437,
	x_18 => x_438,
	x_19 => x_439,
	x_20 => x_440,
	x_21 => x_441,
	x_22 => x_442,
	x_23 => x_443,
	x_24 => x_444,
	x_25 => x_445,
	x_26 => x_446,
	x_27 => x_447,
	y_0 => y_420,
	y_1 => y_421,
	y_2 => y_422,
	y_3 => y_423,
	y_4 => y_424,
	y_5 => y_425,
	y_6 => y_426,
	y_7 => y_427,
	y_8 => y_428,
	y_9 => y_429,
	y_10 => y_430,
	y_11 => y_431,
	y_12 => y_432,
	y_13 => y_433,
	y_14 => y_434,
	y_15 => y_435,
	y_16 => y_436,
	y_17 => y_437,
	y_18 => y_438,
	y_19 => y_439,
	y_20 => y_440,
	y_21 => y_441,
	y_22 => y_442,
	y_23 => y_443,
	y_24 => y_444,
	y_25 => y_445,
	y_26 => y_446,
	y_27 => y_447
    );
ut16_lstm_layer_16: lstm_layer_16 port map(
	x_0 => x_448,
	x_1 => x_449,
	x_2 => x_450,
	x_3 => x_451,
	x_4 => x_452,
	x_5 => x_453,
	x_6 => x_454,
	x_7 => x_455,
	x_8 => x_456,
	x_9 => x_457,
	x_10 => x_458,
	x_11 => x_459,
	x_12 => x_460,
	x_13 => x_461,
	x_14 => x_462,
	x_15 => x_463,
	x_16 => x_464,
	x_17 => x_465,
	x_18 => x_466,
	x_19 => x_467,
	x_20 => x_468,
	x_21 => x_469,
	x_22 => x_470,
	x_23 => x_471,
	x_24 => x_472,
	x_25 => x_473,
	x_26 => x_474,
	x_27 => x_475,
	y_0 => y_448,
	y_1 => y_449,
	y_2 => y_450,
	y_3 => y_451,
	y_4 => y_452,
	y_5 => y_453,
	y_6 => y_454,
	y_7 => y_455,
	y_8 => y_456,
	y_9 => y_457,
	y_10 => y_458,
	y_11 => y_459,
	y_12 => y_460,
	y_13 => y_461,
	y_14 => y_462,
	y_15 => y_463,
	y_16 => y_464,
	y_17 => y_465,
	y_18 => y_466,
	y_19 => y_467,
	y_20 => y_468,
	y_21 => y_469,
	y_22 => y_470,
	y_23 => y_471,
	y_24 => y_472,
	y_25 => y_473,
	y_26 => y_474,
	y_27 => y_475
    );
ut17_lstm_layer_17: lstm_layer_17 port map(
	x_0 => x_476,
	x_1 => x_477,
	x_2 => x_478,
	x_3 => x_479,
	x_4 => x_480,
	x_5 => x_481,
	x_6 => x_482,
	x_7 => x_483,
	x_8 => x_484,
	x_9 => x_485,
	x_10 => x_486,
	x_11 => x_487,
	x_12 => x_488,
	x_13 => x_489,
	x_14 => x_490,
	x_15 => x_491,
	x_16 => x_492,
	x_17 => x_493,
	x_18 => x_494,
	x_19 => x_495,
	x_20 => x_496,
	x_21 => x_497,
	x_22 => x_498,
	x_23 => x_499,
	x_24 => x_500,
	x_25 => x_501,
	x_26 => x_502,
	x_27 => x_503,
	y_0 => y_476,
	y_1 => y_477,
	y_2 => y_478,
	y_3 => y_479,
	y_4 => y_480,
	y_5 => y_481,
	y_6 => y_482,
	y_7 => y_483,
	y_8 => y_484,
	y_9 => y_485,
	y_10 => y_486,
	y_11 => y_487,
	y_12 => y_488,
	y_13 => y_489,
	y_14 => y_490,
	y_15 => y_491,
	y_16 => y_492,
	y_17 => y_493,
	y_18 => y_494,
	y_19 => y_495,
	y_20 => y_496,
	y_21 => y_497,
	y_22 => y_498,
	y_23 => y_499,
	y_24 => y_500,
	y_25 => y_501,
	y_26 => y_502,
	y_27 => y_503
    );
ut18_lstm_layer_18: lstm_layer_18 port map(
	x_0 => x_504,
	x_1 => x_505,
	x_2 => x_506,
	x_3 => x_507,
	x_4 => x_508,
	x_5 => x_509,
	x_6 => x_510,
	x_7 => x_511,
	x_8 => x_512,
	x_9 => x_513,
	x_10 => x_514,
	x_11 => x_515,
	x_12 => x_516,
	x_13 => x_517,
	x_14 => x_518,
	x_15 => x_519,
	x_16 => x_520,
	x_17 => x_521,
	x_18 => x_522,
	x_19 => x_523,
	x_20 => x_524,
	x_21 => x_525,
	x_22 => x_526,
	x_23 => x_527,
	x_24 => x_528,
	x_25 => x_529,
	x_26 => x_530,
	x_27 => x_531,
	y_0 => y_504,
	y_1 => y_505,
	y_2 => y_506,
	y_3 => y_507,
	y_4 => y_508,
	y_5 => y_509,
	y_6 => y_510,
	y_7 => y_511,
	y_8 => y_512,
	y_9 => y_513,
	y_10 => y_514,
	y_11 => y_515,
	y_12 => y_516,
	y_13 => y_517,
	y_14 => y_518,
	y_15 => y_519,
	y_16 => y_520,
	y_17 => y_521,
	y_18 => y_522,
	y_19 => y_523,
	y_20 => y_524,
	y_21 => y_525,
	y_22 => y_526,
	y_23 => y_527,
	y_24 => y_528,
	y_25 => y_529,
	y_26 => y_530,
	y_27 => y_531
    );
ut19_lstm_layer_19: lstm_layer_19 port map(
	x_0 => x_532,
	x_1 => x_533,
	x_2 => x_534,
	x_3 => x_535,
	x_4 => x_536,
	x_5 => x_537,
	x_6 => x_538,
	x_7 => x_539,
	x_8 => x_540,
	x_9 => x_541,
	x_10 => x_542,
	x_11 => x_543,
	x_12 => x_544,
	x_13 => x_545,
	x_14 => x_546,
	x_15 => x_547,
	x_16 => x_548,
	x_17 => x_549,
	x_18 => x_550,
	x_19 => x_551,
	x_20 => x_552,
	x_21 => x_553,
	x_22 => x_554,
	x_23 => x_555,
	x_24 => x_556,
	x_25 => x_557,
	x_26 => x_558,
	x_27 => x_559,
	y_0 => y_532,
	y_1 => y_533,
	y_2 => y_534,
	y_3 => y_535,
	y_4 => y_536,
	y_5 => y_537,
	y_6 => y_538,
	y_7 => y_539,
	y_8 => y_540,
	y_9 => y_541,
	y_10 => y_542,
	y_11 => y_543,
	y_12 => y_544,
	y_13 => y_545,
	y_14 => y_546,
	y_15 => y_547,
	y_16 => y_548,
	y_17 => y_549,
	y_18 => y_550,
	y_19 => y_551,
	y_20 => y_552,
	y_21 => y_553,
	y_22 => y_554,
	y_23 => y_555,
	y_24 => y_556,
	y_25 => y_557,
	y_26 => y_558,
	y_27 => y_559
    );
ut20_lstm_layer_20: lstm_layer_20 port map(
	x_0 => x_560,
	x_1 => x_561,
	x_2 => x_562,
	x_3 => x_563,
	x_4 => x_564,
	x_5 => x_565,
	x_6 => x_566,
	x_7 => x_567,
	x_8 => x_568,
	x_9 => x_569,
	x_10 => x_570,
	x_11 => x_571,
	x_12 => x_572,
	x_13 => x_573,
	x_14 => x_574,
	x_15 => x_575,
	x_16 => x_576,
	x_17 => x_577,
	x_18 => x_578,
	x_19 => x_579,
	x_20 => x_580,
	x_21 => x_581,
	x_22 => x_582,
	x_23 => x_583,
	x_24 => x_584,
	x_25 => x_585,
	x_26 => x_586,
	x_27 => x_587,
	y_0 => y_560,
	y_1 => y_561,
	y_2 => y_562,
	y_3 => y_563,
	y_4 => y_564,
	y_5 => y_565,
	y_6 => y_566,
	y_7 => y_567,
	y_8 => y_568,
	y_9 => y_569,
	y_10 => y_570,
	y_11 => y_571,
	y_12 => y_572,
	y_13 => y_573,
	y_14 => y_574,
	y_15 => y_575,
	y_16 => y_576,
	y_17 => y_577,
	y_18 => y_578,
	y_19 => y_579,
	y_20 => y_580,
	y_21 => y_581,
	y_22 => y_582,
	y_23 => y_583,
	y_24 => y_584,
	y_25 => y_585,
	y_26 => y_586,
	y_27 => y_587
    );
ut21_lstm_layer_21: lstm_layer_21 port map(
	x_0 => x_588,
	x_1 => x_589,
	x_2 => x_590,
	x_3 => x_591,
	x_4 => x_592,
	x_5 => x_593,
	x_6 => x_594,
	x_7 => x_595,
	x_8 => x_596,
	x_9 => x_597,
	x_10 => x_598,
	x_11 => x_599,
	x_12 => x_600,
	x_13 => x_601,
	x_14 => x_602,
	x_15 => x_603,
	x_16 => x_604,
	x_17 => x_605,
	x_18 => x_606,
	x_19 => x_607,
	x_20 => x_608,
	x_21 => x_609,
	x_22 => x_610,
	x_23 => x_611,
	x_24 => x_612,
	x_25 => x_613,
	x_26 => x_614,
	x_27 => x_615,
	y_0 => y_588,
	y_1 => y_589,
	y_2 => y_590,
	y_3 => y_591,
	y_4 => y_592,
	y_5 => y_593,
	y_6 => y_594,
	y_7 => y_595,
	y_8 => y_596,
	y_9 => y_597,
	y_10 => y_598,
	y_11 => y_599,
	y_12 => y_600,
	y_13 => y_601,
	y_14 => y_602,
	y_15 => y_603,
	y_16 => y_604,
	y_17 => y_605,
	y_18 => y_606,
	y_19 => y_607,
	y_20 => y_608,
	y_21 => y_609,
	y_22 => y_610,
	y_23 => y_611,
	y_24 => y_612,
	y_25 => y_613,
	y_26 => y_614,
	y_27 => y_615
    );
ut22_lstm_layer_22: lstm_layer_22 port map(
	x_0 => x_616,
	x_1 => x_617,
	x_2 => x_618,
	x_3 => x_619,
	x_4 => x_620,
	x_5 => x_621,
	x_6 => x_622,
	x_7 => x_623,
	x_8 => x_624,
	x_9 => x_625,
	x_10 => x_626,
	x_11 => x_627,
	x_12 => x_628,
	x_13 => x_629,
	x_14 => x_630,
	x_15 => x_631,
	x_16 => x_632,
	x_17 => x_633,
	x_18 => x_634,
	x_19 => x_635,
	x_20 => x_636,
	x_21 => x_637,
	x_22 => x_638,
	x_23 => x_639,
	x_24 => x_640,
	x_25 => x_641,
	x_26 => x_642,
	x_27 => x_643,
	y_0 => y_616,
	y_1 => y_617,
	y_2 => y_618,
	y_3 => y_619,
	y_4 => y_620,
	y_5 => y_621,
	y_6 => y_622,
	y_7 => y_623,
	y_8 => y_624,
	y_9 => y_625,
	y_10 => y_626,
	y_11 => y_627,
	y_12 => y_628,
	y_13 => y_629,
	y_14 => y_630,
	y_15 => y_631,
	y_16 => y_632,
	y_17 => y_633,
	y_18 => y_634,
	y_19 => y_635,
	y_20 => y_636,
	y_21 => y_637,
	y_22 => y_638,
	y_23 => y_639,
	y_24 => y_640,
	y_25 => y_641,
	y_26 => y_642,
	y_27 => y_643
    );
ut23_lstm_layer_23: lstm_layer_23 port map(
	x_0 => x_644,
	x_1 => x_645,
	x_2 => x_646,
	x_3 => x_647,
	x_4 => x_648,
	x_5 => x_649,
	x_6 => x_650,
	x_7 => x_651,
	x_8 => x_652,
	x_9 => x_653,
	x_10 => x_654,
	x_11 => x_655,
	x_12 => x_656,
	x_13 => x_657,
	x_14 => x_658,
	x_15 => x_659,
	x_16 => x_660,
	x_17 => x_661,
	x_18 => x_662,
	x_19 => x_663,
	x_20 => x_664,
	x_21 => x_665,
	x_22 => x_666,
	x_23 => x_667,
	x_24 => x_668,
	x_25 => x_669,
	x_26 => x_670,
	x_27 => x_671,
	y_0 => y_644,
	y_1 => y_645,
	y_2 => y_646,
	y_3 => y_647,
	y_4 => y_648,
	y_5 => y_649,
	y_6 => y_650,
	y_7 => y_651,
	y_8 => y_652,
	y_9 => y_653,
	y_10 => y_654,
	y_11 => y_655,
	y_12 => y_656,
	y_13 => y_657,
	y_14 => y_658,
	y_15 => y_659,
	y_16 => y_660,
	y_17 => y_661,
	y_18 => y_662,
	y_19 => y_663,
	y_20 => y_664,
	y_21 => y_665,
	y_22 => y_666,
	y_23 => y_667,
	y_24 => y_668,
	y_25 => y_669,
	y_26 => y_670,
	y_27 => y_671
    );
ut24_lstm_layer_24: lstm_layer_24 port map(
	x_0 => x_672,
	x_1 => x_673,
	x_2 => x_674,
	x_3 => x_675,
	x_4 => x_676,
	x_5 => x_677,
	x_6 => x_678,
	x_7 => x_679,
	x_8 => x_680,
	x_9 => x_681,
	x_10 => x_682,
	x_11 => x_683,
	x_12 => x_684,
	x_13 => x_685,
	x_14 => x_686,
	x_15 => x_687,
	x_16 => x_688,
	x_17 => x_689,
	x_18 => x_690,
	x_19 => x_691,
	x_20 => x_692,
	x_21 => x_693,
	x_22 => x_694,
	x_23 => x_695,
	x_24 => x_696,
	x_25 => x_697,
	x_26 => x_698,
	x_27 => x_699,
	y_0 => y_672,
	y_1 => y_673,
	y_2 => y_674,
	y_3 => y_675,
	y_4 => y_676,
	y_5 => y_677,
	y_6 => y_678,
	y_7 => y_679,
	y_8 => y_680,
	y_9 => y_681,
	y_10 => y_682,
	y_11 => y_683,
	y_12 => y_684,
	y_13 => y_685,
	y_14 => y_686,
	y_15 => y_687,
	y_16 => y_688,
	y_17 => y_689,
	y_18 => y_690,
	y_19 => y_691,
	y_20 => y_692,
	y_21 => y_693,
	y_22 => y_694,
	y_23 => y_695,
	y_24 => y_696,
	y_25 => y_697,
	y_26 => y_698,
	y_27 => y_699
    );
ut25_lstm_layer_25: lstm_layer_25 port map(
	x_0 => x_700,
	x_1 => x_701,
	x_2 => x_702,
	x_3 => x_703,
	x_4 => x_704,
	x_5 => x_705,
	x_6 => x_706,
	x_7 => x_707,
	x_8 => x_708,
	x_9 => x_709,
	x_10 => x_710,
	x_11 => x_711,
	x_12 => x_712,
	x_13 => x_713,
	x_14 => x_714,
	x_15 => x_715,
	x_16 => x_716,
	x_17 => x_717,
	x_18 => x_718,
	x_19 => x_719,
	x_20 => x_720,
	x_21 => x_721,
	x_22 => x_722,
	x_23 => x_723,
	x_24 => x_724,
	x_25 => x_725,
	x_26 => x_726,
	x_27 => x_727,
	y_0 => y_700,
	y_1 => y_701,
	y_2 => y_702,
	y_3 => y_703,
	y_4 => y_704,
	y_5 => y_705,
	y_6 => y_706,
	y_7 => y_707,
	y_8 => y_708,
	y_9 => y_709,
	y_10 => y_710,
	y_11 => y_711,
	y_12 => y_712,
	y_13 => y_713,
	y_14 => y_714,
	y_15 => y_715,
	y_16 => y_716,
	y_17 => y_717,
	y_18 => y_718,
	y_19 => y_719,
	y_20 => y_720,
	y_21 => y_721,
	y_22 => y_722,
	y_23 => y_723,
	y_24 => y_724,
	y_25 => y_725,
	y_26 => y_726,
	y_27 => y_727
    );
ut26_lstm_layer_26: lstm_layer_26 port map(
	x_0 => x_728,
	x_1 => x_729,
	x_2 => x_730,
	x_3 => x_731,
	x_4 => x_732,
	x_5 => x_733,
	x_6 => x_734,
	x_7 => x_735,
	x_8 => x_736,
	x_9 => x_737,
	x_10 => x_738,
	x_11 => x_739,
	x_12 => x_740,
	x_13 => x_741,
	x_14 => x_742,
	x_15 => x_743,
	x_16 => x_744,
	x_17 => x_745,
	x_18 => x_746,
	x_19 => x_747,
	x_20 => x_748,
	x_21 => x_749,
	x_22 => x_750,
	x_23 => x_751,
	x_24 => x_752,
	x_25 => x_753,
	x_26 => x_754,
	x_27 => x_755,
	y_0 => y_728,
	y_1 => y_729,
	y_2 => y_730,
	y_3 => y_731,
	y_4 => y_732,
	y_5 => y_733,
	y_6 => y_734,
	y_7 => y_735,
	y_8 => y_736,
	y_9 => y_737,
	y_10 => y_738,
	y_11 => y_739,
	y_12 => y_740,
	y_13 => y_741,
	y_14 => y_742,
	y_15 => y_743,
	y_16 => y_744,
	y_17 => y_745,
	y_18 => y_746,
	y_19 => y_747,
	y_20 => y_748,
	y_21 => y_749,
	y_22 => y_750,
	y_23 => y_751,
	y_24 => y_752,
	y_25 => y_753,
	y_26 => y_754,
	y_27 => y_755
    );
        y_0 <= "0000000000000000";

        y_1 <= "0000000000000000";

        y_2 <= "0000000000000000";

        y_3 <= "0000000000000000";

        y_4 <= "0000000000000000";

        y_5 <= "0000000000000000";

        y_6 <= "0000000000000000";

        y_7 <= "0000000000000000";

        y_8 <= "0000000000000000";

        y_9 <= "0000000000000000";

        y_10 <= "0000000000000000";

        y_11 <= "0000000000000000";

        y_12 <= "0000000000000000";

        y_13 <= "0000000000000000";

        y_14 <= "0000000000000000";

        y_15 <= "0000000000000000";

        y_16 <= "0000000000000000";

        y_17 <= "0000000000000000";

        y_18 <= "0000000000000000";

        y_19 <= "0000000000000000";

        y_20 <= "0000000000000000";

        y_21 <= "0000000000000000";

        y_22 <= "0000000000000000";

        y_23 <= "0000000000000000";

        y_24 <= "0000000000000000";

        y_25 <= "0000000000000000";

        y_26 <= "0000000000000000";

        y_27 <= "0000000000000000";

        y_28 <= "0000000000000000";

        y_29 <= "0000000000000000";

        y_30 <= "0000000000000000";

        y_31 <= "0000000000000000";

        y_32 <= "0000000000000000";

        y_33 <= "0000000000000000";

        y_34 <= "0000000000000000";

        y_35 <= "0000000000000000";

        y_36 <= "0000000000000000";

        y_37 <= "0000000000000000";

        y_38 <= "0000000000000000";

        y_39 <= "0000000000000000";

        y_40 <= "0000000000000000";

        y_41 <= "0000000000000000";

        y_42 <= "0000000000000000";

        y_43 <= "0000000000000000";

        y_44 <= "0000000000000000";

        y_45 <= "0000000000000000";

        y_46 <= "0000000000000000";

        y_47 <= "0000000000000000";

        y_48 <= "0000000000000000";

        y_49 <= "0000000000000000";

        y_50 <= "0000000000000000";

        y_51 <= "0000000000000000";

        y_52 <= "0000000000000000";

        y_53 <= "0000000000000000";

        y_54 <= "0000000000000000";

        y_55 <= "0000000000000000";

        y_56 <= "0000000000000000";

        y_57 <= "0000000000000000";

        y_58 <= "0000000000000000";

        y_59 <= "0000000000000000";

        y_60 <= "0000000000000000";

        y_61 <= "0000000000000000";

        y_62 <= "0000000000000000";

        y_63 <= "0000000000000000";

        y_64 <= "0000000000000000";

        y_65 <= "0000000000000000";

        y_66 <= "0000000000000000";

        y_67 <= "0000000000000000";

        y_68 <= "0000000000000000";

        y_69 <= "0000000000000000";

        y_70 <= "0000000000000000";

        y_71 <= "0000000000000000";

        y_72 <= "0000000000000000";

        y_73 <= "0000000000000000";

        y_74 <= "0000000000000000";

        y_75 <= "0000000000000000";

        y_76 <= "0000000000000000";

        y_77 <= "0000000000000000";

        y_78 <= "0000000000000000";

        y_79 <= "0000000000000000";

        y_80 <= "0000000000000000";

        y_81 <= "0000000000000000";

        y_82 <= "0000000000000000";

        y_83 <= "0000000000000000";

        y_84 <= "0000000000000000";

        y_85 <= "0000000000000000";

        y_86 <= "0000000000000000";

        y_87 <= "0000000000000000";

        y_88 <= "0000000000000000";

        y_89 <= "0000000000000000";

        y_90 <= "0000000000000000";

        y_91 <= "0000000000000000";

        y_92 <= "0000000000000000";

        y_93 <= "0000000000000000";

        y_94 <= "0000000000000000";

        y_95 <= "0000000000000000";

        y_96 <= "0000000000000000";

        y_97 <= "0000000000000000";

        y_98 <= "0000000000000000";

        y_99 <= "0000000000000000";

        y_100 <= "0000000000000000";

        y_101 <= "0000000000000000";

        y_102 <= "0000000000000000";

        y_103 <= "0000000000000000";

        y_104 <= "0000000000000000";

        y_105 <= "0000000000000000";

        y_106 <= "0000000000000000";

        y_107 <= "0000000000000000";

        y_108 <= "0000000000000000";

        y_109 <= "0000000000000000";

        y_110 <= "0000000000000000";

        y_111 <= "0000000000000000";

        y_756 <= "0000000000000000";

        y_757 <= "0000000000000000";

        y_758 <= "0000000000000000";

        y_759 <= "0000000000000000";

        y_760 <= "0000000000000000";

        y_761 <= "0000000000000000";

        y_762 <= "0000000000000000";

        y_763 <= "0000000000000000";

        y_764 <= "0000000000000000";

        y_765 <= "0000000000000000";

        y_766 <= "0000000000000000";

        y_767 <= "0000000000000000";

        y_768 <= "0000000000000000";

        y_769 <= "0000000000000000";

        y_770 <= "0000000000000000";

        y_771 <= "0000000000000000";

        y_772 <= "0000000000000000";

        y_773 <= "0000000000000000";

        y_774 <= "0000000000000000";

        y_775 <= "0000000000000000";

        y_776 <= "0000000000000000";

        y_777 <= "0000000000000000";

        y_778 <= "0000000000000000";

        y_779 <= "0000000000000000";

        y_780 <= "0000000000000000";

        y_781 <= "0000000000000000";

        y_782 <= "0000000000000000";

        y_783 <= "0000000000000000";
end Behavioral;