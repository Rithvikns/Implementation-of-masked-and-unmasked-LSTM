library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_2 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_2;

architecture syn of ram_2 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"0000000000011011","0000000010111011","0000000000100001","0000000011110000","0000000010011110","0000000111111000","0000000111111111","0000000101101110","1000000111000101","0000000011110100","1000000111110011","1000000000101101","1000100011000001","1000010110111110","0000101010100110","0000001010010011","1000000101110110","1000000110001100","1000000110111010","1000000001000010","1000000001011110","1000000001001011","0000000111011010","1000000001110000","0000000001101101","1000000111011100","0000000010101101","1000000000101110","0000000111100001","0000000011101101","1000000000111011","0000000011010010","1000011100101000","1000101011010011","1001101000100010","1001111111000100","1001000101100111","1000111101010001","1000110010000001","1001001010010000","1001111110011011","1001001100100011","1000100100000111","0000001110100100","0001011100100000","1000000111100110","1001011110001001","1001100101110111","1010011011001010","1001100100001110","1000111000111111","1000011111101101","0000000000101011","0000000010100001","1000000000111101","1000000011010011","1000000010000110","0000000000010100","1000010111000000","1000101000111100","1001010001011101","0000011010100010","0000100001010010","1001011100011000","0000100101000110","0000101010111100","0000001111000110","0000011001001010","0000101011011001","1000000011100010","1000100001001000","1000000001100111","1000000000100110","1000001101000010","1000100100010001","1001010101110100","1000111110010100","1000100011010100","1010010111010101","0000001101001111","0000111001110100","0000101110100010","1000000101110111","1000000011011110","1000000000111001","0000000100111000","0000000110000100","1001001110011010","1000101101010000","0000000000000110","0000001001100111","1000011100110000","0000011111000100","0001001001111101","0000000101101000","0000011110010001","0000100001111110","0000110110101001","0000011110110110","0000000010101011","1000000001000010","1000000011110001","1000100111001001","1000110101011010","1000111101011101","1000101000001101","1000000100001011","1000101000010100","1000011010001110","0000010000101101","1000110000111100","1000000001001100","0000000000001001","1000101101100111","1000100110011111","1000111100111101","1000101011001111","0000001010110010","0000101110111011","0000001000001100","0000010110100101","0000110110101010","0000000110110100","0000000101011101","0000010101001011","0000001001110100","0000010000111011","1000001000010000","0000000011100010","0000000101100110","1000001001111011","1000100111100100","1000101111000001","1000100110011000","1001000000101001","1001000001001001","1010000010001000","0000010111110001","1001010000000010","1000101101111010","1000000010111010","1000000100110001","0000011110001111","0000011100100011","1000000001011001","1000000001101001","1000010000011111","1000000101010011","1000000111101001","0000001010000101","0000011000001110","0000000000010011","1000001101011110","1000001011100010","1000001011110000","1000000100100101","0000010010000100","1000000011000010","1000000000110101","1000010111000111","1000010111010110","0000001000110000","1000001000111001","1000001000011010","1001001000001011","0000001110101111","1001110111011001","1000111010111010","0000000101101011","1000100101111011","1000101101101101","1000000010010011","0000000011010100","1000001101011010","0000000010100010","0000000101011011","1000000101100100","0000001011100111","0000001101001110","1000010000100101","1000011001001011","1000011011110101","1000010001011010","1000001001100101","1000001011110000","1000010110101010","1000010101011011","1000011100101101","1000011100010010","1000100100001101","1000010100101111","1000110000101011","1001001000001101","1001001000101001","1000011100011001","1000101101011111","0000000001110110","1001101001010101","0000010011111110","0000000010101110","0000001111010101","0000000111110001","0000000010111100","0000000001110001","0000001101001100","1000001100010010","1000000100111101","0000001111010111","1000100011001100","1000001000101011","1000011010010001","1000100101001100","1000100001110100","1000111010100011","1000100110010010","1000010011001101","1000101100011011","0000010011100010","0000011011000110","1000110101110100","1001011101101001","1001011110000111","1000101111100010","1000111000100001","1000110010111011","0000101110011101","0000000010111101","1000001111010010","0000010101000001","1000001010111110","1000011001001110","1000001101110011","1000010011010011","1000010101110001","0000011010010010","1000001111100110","1000100000000110","1000100111111110","1000101001100011","1000100100111110","1000111010010000","1000010011011110","1000111010010001","1000000110000000","1000000100011111","1000001100110101","1000011100101111","1000010000100010","1000111000111101","1010101110011011","1001011000000111","1000101000101001","0000000010000110","1001011010000100","1000110011111000","1000000001001110","0000001101100011","0000001100010000","1000010110110011","1000010110001001","1000010001000010","1000001011011001","0000000011101010","1000001111011101","1000011101000011","1000110000000010","1000011000101011","1000001111000001","1000011010111011","1000010010101100","1000011111100111","1000010010110011","0000000100001111","1000101111101111","1000001101101010","1000010001110101","1001011101000111","1001111000010110","1000010011101010","1001000111101011","1000000000110001","1001000010101100","1000101011011000","0000011010100010","1000010011010101","0000100011010110","0000101011000101","1000011100110110","1000001111000001","1000011111010100","1000011111011111","1000000011001101","1000010011101001","1000110011100110","1000011101000001","1000110111110111","1000010111100101","0000001011111101","1000010100010101","1000010001000011","1000000010110010","1000011101111100","1000011100101111","1000110001011110","1001011000111110","1000001010101010","0000010010000101","1001010000111010","1000000110001100","1001010011111111","1001011101100011","1000110000110100","1000011000110010","0000100011100110","0000001011010001","1001001101010011","1001000000101100","1001101111001111","1010001001001011","1001101110010101","1001111011101010","1010111000110111","1010001111100110","1001100010101110","1000110000100111","1000110100110000","1000100100101110","0000001011011000","1000010000010001","0000000110010011","1000001001011110","1000001111111101","1000101111010010","0000011110010110","1001001010000111","1000111100010101","1000000101111000","1001000000111010","1001110101010010","1001101011100000","1000010110010011","1000111110000010","1010010000110011","1010100100101100","1001111111100000","1001111101101110","1001101110011100","1001100111001111","1001101111010100","1001111000100100","1010000000011011","1001110111001010","1001001101111101","1000111000110000","1000111001001100","0000000010110111","1000001111100010","0000000110110010","1000100101100000","1000111010010000","0000011110001011","0000111101111001","0000101111000111","1000001100111011","1000100100011110","1000111010010100","0000000101001100","1001001010100110","1010101010010001","1011000011010110","1011011010111100","1010000101001000","1001001010101010","1000101000111000","1000011010100101","0000010011101101","1000000101100101","1000010100000001","1000101100000110","1001011101100010","1001000000111010","1000101000110110","1000101111001001","1000010100011111","1000011001111111","1000011000111010","1000010000110000","1000001000000010","0001010010011010","0001010000011100","0010001010111111","0000111110111000","1000101110100101","1001010010000001","1000111011111101","1001001001100101","1001110010010010","1001111001111100","1001001101010111","1000010001111111","1000001010100101","1000001001001111","1000000101000011","0000001010100001","1000000010100011","1000000001000010","1000100110010110","1000111010001010","1000111011111010","1000110011100011","1000001101010101","1000110010110101","1000001110010000","1000101111001000","1000000010101101","1000000101001111","0000000110110011","0000011101111010","0001100110110010","0001001010111010","1000011111010111","1000110111000110","1000110101000001","1000001100100011","0000001011101011","0001010110100000","0000011101001111","1000001110101001","1000001110000011","1000000010110001","1000000001010001","1000000111111111","1000010100010001","0000000010101011","1000010011101101","1000101110101101","1000101101101110","1000100101010011","1000100000110001","0000000101000011","1000001000101110","0000000011001111","1000010110110010","1000010010001001","0000101001110010","0001000111011100","0001000110000100","0001011001100101","0000000010111011","1001001000110000","0000000110100110","0000010101110110","0000001000110110","0000101101110011","0000010001101111","1000001111110010","1000010011010000","0000001111001101","0000000100010010","0000001111011100","0000011110101101","0000011101100110","1000001101010011","1000011011100101","1000000010111000","0000010100010111","1000010111010111","1000010010000000","1000010101011000","0000010111000100","0000010011111101","0000100111010001","0000101100101110","0001111001100011","0010000011000000","0001100001100001","0000000001111110","1001001101101011","0000100111100000","0000000100101011","0000001100000010","0000011000111100","0000010110000110","1000000101100001","0000000001111100","0000001100110001","0000100001010100","0000011000110101","0000100111010111","0000000100010101","1000100101000001","1000010100010100","1000011010100001","1000011111100101","1000010001110110","1000100001001101","1000000100101100","0000000110010110","1000001000100110","1000000110110001","1000000011000000","0001000001011111","0000011101011000","0001111110011111","1000101010011011","1001000001011111","1000010011011100","0000000001011010","0000001000100101","0000011100001011","0000010110101000","0000001100111101","0000010011110001","1000001001010101","0000000111101110","1000000010010001","0000100011011111","0000001000110110","1000100000100101","1000101110110011","1000010011110000","0000001001101110","0000000010100101","1000000111011001","1000001011010011","1000000001010001","0000011000001011","0000011100111110","0001000100011001","0000011111101011","1000110101000111","0000110011011100","1000110000100001","1001000001100101","1000111110011110","1000100000010000","0000000001000000","1000010001101001","0000000111010100","0000010000001100","0000010011011010","0000001100011111","0000011010001110","0000001100110000","0000001111111001","0000001110010110","1000001110011001","1000000100100100","0000001011000110","0000011001000010","0000000011101011","1000010111010010","1000001000111101","0000000110001101","0000101011000010","1000001001000000","0000010001001111","0000101111011111","0001010111110001","0000001010011111","0000000000101000","1000110110100101","1000001001000001","1000000000101001","0000011111011101","0000001001101010","0000100100110101","0000000110011101","0000100000100100","0000001010011100","0000010101110000","0000101101110110","0000001001000110","1000010010100011","1000010010001000","1000001111000010","1000010111001000","1000011111101011","0000001001110010","0000001100010011","0000100111000010","0000010111000010","0000011101111100","0000011011000010","0000011110101000","0000000011001010","0000011110110001","1000110100101101","1000101001111110","0000001011010001","1000001101101010","1000001101111010","1000000010010101","1000001101001111","0000001110111100","1000001001101111","1000000000110010","0000010000110001","0000000101010100","0000001000100000","1000001101010001","1000010010001101","1000010001110111","1000101110101000","1000011010111001","0000001010101101","0000011111000010","0000111010100100","0000001101011110","0000010101000010","0000010010101011","0001011110111110","0000010001010000","1000001001100011","0000001110001000","1000011001011011","1000101101100110","1000101111001011","0000101101110101","0000000011101111","0000010101000011","0000001011100000","0000010100111111","0000001110111110","0000001101001000","0000011001010001","1000000100101100","0000000100011000","0000001110011111","1000010111111110","1000101000110101","1000110101011110","1000100101010001","1000010010011111","0000011001111111","0000001111110111","0000001111101110","0000010000100111","0000110110101111","0000000101100111","0000100001011000","0000001000010010","1000111010111010","1000100111111000","0000000110100111","0000000010000101","1000101101110101","1000110110111101","1000010110111001","0000111000101110","0000010000111111","0000000111110101","1000000011111111","0000000001101100","1000011010111001","0000000011100101","0000001000100100","1000100010010010","1000100111101000","1000110001011011","1000101011110010","1000010111111101","0000011111010101","0000100101111100","0000011111010010","0000100110110011","0001001000000101","0000010000010010","0000100010011101","0000100110011111","1000111000100110","0000000000111001","0000000000100011","1000000011100100","1001000001101100","1001110101100111","1000111101101101","1001010111001011","1000110011011010","1000110001010011","1000001111111111","1000101011001011","1000100010010101","0000000100011000","0000101000011000","1000010011001011","0000010010001011","1000010111101000","1000100011110101","1000010111100001","0000010101011110","0000101000111100","0000011010001100","0000101011110001","0000000110110001","1000101011111110","0000101110001111","0001111001111001","0000100001110100","1000000000110000","1000000111101000","1000000110000010","1000100101100111","1001000110100110","1010100001011100","1010110000100101","1000110101001010","1001001111011010","1010101010111111","1011001111101011","1010010010100011","1001111101001010","1001100010000100","1001001101111011","1000011011001010","1000000000110111","1000000100001110","1000010111011000","1000111000010001","1001100110010110","1000100110110101","0000001110110101","1000100000001001","1010000100010001","1010010111100001","0000110001001111","0000101100111011","1000000111100110","0000000011101010","0000000011101001","0000000011011111","1000001100011011","1001011011000100","1001011010000111","1001011000101010","1001110010100101","1001111111000111","1001111000010110","1010111011100110","1001100010110000","1011100110000100","1011100110011011","1011111000011000","1010111111000101","1010110011110110","1010010000100001","1010101000101111","1001110000011101","1001101001010000","1001101011001100","1001110111101101","1000111110001100","1000001011110100","1000001100111111","0000000010110101","0000000011010100","0000000111101101","0000000001000000","0000000011111110","0000000001010110","1000000011111111","1000001000000000","1000001010110100","1000011011011101","1000011111110011","1000101000000101","1001000001001101","1001010111000111","1000111101101000","1001001100101010","1001001110001000","1001001000101101","1001000011111001","1001010000111110","1001011110111011","1000101000011100","1000111111111100","1001001001111010","1000111011000101","1000001101000000","1000000110010101","1000000010101100","0000000001010010","1000000011110001");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
