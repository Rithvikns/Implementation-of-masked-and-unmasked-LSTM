library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_1 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_1;

architecture syn of ram_1 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"0000000110000101","1000000000100010","0000000110001111","0000000010011001","1000000011101101","1000000100011011","1000000100111100","0000000111001010","0000000100000010","1000000011011100","0000000000101100","1000000110011111","1000000110011001","1000010100110010","1000000011100101","0000000011100010","1000000001001110","0000000100101000","1000000001111010","0000000011100100","1000000110011001","0000000010000001","1000000000101110","0000000100101111","0000000000010101","0000000010000011","1000000000110001","0000000110110001","0000000101011001","0000000100100111","0000000010011011","1000000110000010","0000000010101010","0000000011101111","0000000010100011","1000011110111001","1000110000111101","1000111010010001","1001011011111100","1001001010111111","1001000110110101","1001101001101100","0001000010111111","0000101101110001","1000111101100001","1001101101000000","1000111100110011","1000011111001000","1000010100100010","1000000111100001","0000000011001101","0000000010110100","1000000000011000","1000000001101010","0000000010100111","1000000001000101","0000000111111100","1000000001000011","0000000001010001","1000000000010010","1000001100010111","1000100110101001","1000101100101101","1001100010101011","1001000100101000","1001011011000100","1001100111111111","1010110101101111","1001000100111011","0000101101110110","0001010010011101","0001100110100111","0001011111111110","1000011000100011","1000111000100001","1000011111001111","1000010011010100","1010001111110011","1001001101101100","1000111000011110","1000111101011101","1000011100000001","0000000010110011","0000000000100110","1000000100100110","1000000011101011","0000110011101000","0000110000101001","1000110010010000","1001010101111000","1010001101001010","1001000001001001","1010000010011000","1001001001101010","1001110110100011","1010011001010110","1001000101001111","0000000101110101","1000011011010001","1000000110001100","0000010010011010","1001100100100100","1001100000000001","1000111000011000","1000110101101110","1001000100001100","1000110100110011","1001101010101101","1010011100100001","1001001000000010","1000110001001010","0000000110111010","0000000001011100","1000000011001011","0000101100100110","1000000001000100","0000100000100110","1000010000111011","1000101010001111","1000001110110100","0000000010111011","1000011100110101","1000010000101110","1000110100011001","1001000001101101","1000010100000011","1000010000011001","1000010010011100","1000001110011100","1000101110011011","1000110100011111","1000001110101011","1000001110110001","1000001101100011","1000101010100110","1000010100111110","1000101111001111","1010010000001110","1001100011111001","1000110101000010","1000000010100110","0000000011101100","0001000100100100","0000110111011001","0001001110000010","0000011001110011","0000011100010011","1000010001001010","1000110101100110","1000110110111011","1001010001111001","1001011100000100","1001011101101001","1000101110011110","1000111101011011","1000000010000111","1000010111101000","1001001000100001","1001001001001101","1000101100010101","1000100011010110","0000001010111101","0000000100010110","1000011000111111","0000000010000111","1001000110111010","1000110010101010","1000110101000111","1000000000101011","1000010011100100","1001010011110110","1000001101101011","0001100110000111","1000101110000000","1000000001001000","1001001011000010","1001000001011110","1000111111110111","1000110011110000","1000010000100100","1000111100100001","1000111101101001","1001001100100101","1001000101010000","1000111110010001","1001000100001111","1000101111100111","1000011110110000","1000011110010001","1000001101101001","1000011100010111","1000011011001100","1000000011001101","1010111001110110","1001101000110011","1000100010011111","0000000011001000","1000111100011101","1000110000011101","1000100100010000","0000001101000100","1001001111010000","1001011000100111","1000101011011100","1001011001111011","1000001110011101","1000111010111011","1000111010010100","1000100010110100","1001000110000101","1000010111001010","1001000111111001","1000111101010111","1000110101001111","1001001011110011","1000010011001010","1000010110100010","0000000100000011","1000011000100000","1000001111101000","1001000101011100","1001111100100010","0000000001000001","1000100100100110","1000010100100111","1000110110010110","1000110011000111","0000000110010000","1000011111000000","1001001001011011","1000000100111101","1001000001110000","1001001001100001","1000110000010111","1000100100011110","1001001110110111","1000110011101101","1000100010111011","0000001000101110","1000000010100001","1001001111010000","1000110000000010","1000111001000100","1000011100011010","1000101010011101","1000110111000100","1000010000101000","1000101000011000","1010000110011101","1011101000010110","1010011011001010","1000100000110010","1000010110100001","1000110110001010","1000111100000001","1001000000111100","1001000000101100","1000101101111111","1000000100101011","1000100110110001","1001000011000110","1001001010111000","1001001010100110","1001000001000000","1000111010001100","1000001100111100","0000110111000000","0001000001010001","1000001110101101","1001000111001001","1000111110001001","1000110101100000","1000110101100111","1000011100100010","1000101001110100","1000110010111111","1000100100001010","1011000111111011","0000010001110101","1000111001101001","1000010111001111","1000010011101011","1000111000100111","1001010001010101","1000101110000111","1000110101110011","1001010001100101","1000110010010111","1000101101110000","1001000001101001","1000111101011010","1000100010001010","1000101001000000","0000011100101001","0001100001010011","0001110000100111","0000001111101100","1000101010110100","1001001010111101","1000111011110110","1000101011000001","1000001100111101","1000000101111010","1000111100100101","1100111001100111","0000000010110110","0000100011100101","0000110011101100","1000000000011010","0000100111001101","0001000100101111","1001000011100010","1000000101011000","1000000111001011","1010000000110100","1000100010111001","1000101000101001","1000101011100001","1000101001101100","1000101000110000","1000100101111011","0000101000001100","0001101100110011","0001110110011011","0000001110000001","1000101010100010","1000100001110000","1000110001101000","1000101100100111","1001000101010110","1000000100100110","1000101011000101","1001110011011111","1000010011110100","0000101010010111","0000110011111100","0000000011011110","1001000001000110","1000110110000101","0000000111110011","0000001001111010","1000100011011110","1001000110010001","1000110111000111","1000001110010110","1000011110110001","1001100000000001","1001000111110111","1000011110010101","0000100010110001","0010000010110011","0001011111111111","1000000010111010","1000010100011111","1000100011001010","1001100011111001","1000010101000111","1000001010011110","0000101101100011","1000001001000110","1001010101100110","1000100000000000","1000011100100001","1000010001111110","0000101001110100","1000101011101001","1000110111000111","0000101101100111","1000010111010111","1000110101011000","1000111001001100","1000101010011001","0000000000100000","1000000100101001","1001100000110010","1001010111010111","1000010110101110","0000100111111100","0001010100001011","0001001000010100","0000010000001011","0000000100011011","1001101110011000","1001100010011110","0000000000101111","1001010011010010","1000101101010100","1001110000000100","1001100010011100","1000100010100000","1000010101101001","1000111000101101","1000101001101010","1000010101011100","0000101110110001","0001001010111000","0001001101101011","1001001110001000","1000111001000100","1000010100101100","0000010011000101","1001001010011101","1001110011010000","1001101011110111","1000011011111111","0000101111100111","0001010011011010","0001000001011101","0000010100100001","1000101100010000","1001010110100001","1000110011101001","0000000001001111","1000011100111100","0000011111011000","1000010011111111","1000001110101111","0000110011000010","0000100100101001","1000100110000111","1000100110111111","1000000111111110","0000111001111010","0001100101000001","0000110001001110","1001110001110111","1001001100100001","0000011111101011","0000000010111001","1000101010101001","1001110000100110","1000011010010111","0000000101111100","0000110000101010","0001011010001110","0000100010010000","0000011000010110","1001101011011010","1010100011011001","1010001011101000","1001110110001110","1001010100101000","1000101001011011","1001111011000101","1001100010000001","0000100100001111","0000001110110101","1000111001000101","0000000000000000","0000111000010110","0001000100101000","1000101011011011","1000000001011101","1000011100001111","1000001010111100","0000000011000010","1000010010001111","1000011101110001","1000100110000110","1000101000100110","1001000000001100","0000100000011110","0001100010110010","1000000100010100","1000101001010110","1010011111000000","1010010100110011","1001111001110111","1000111010010011","1000110001011010","1000100111000101","1000110101011000","0000001001111001","1010010001111111","1000100110001001","1001010101000101","1000000001000110","0001000001011111","0000100010101011","1001110001011110","1000011110101000","1000100000110001","1000101000101000","1000100110011011","1000101111000001","1000110110101010","1000011111000111","1000111111100110","1000101000100000","0000101001111011","0001100100110011","1000001001001101","1001100000001100","1001101011110110","1001001011001111","0000000111001001","0000001011100001","1000101000110100","0000000110110110","0000010000111111","0000001000110011","1001001111000101","1000101000001010","1001010001111001","1000110111101100","0000110001111111","1001001000110011","1010101111100000","1010001001111111","1001100011010101","1001010100110000","1000101011010110","1000000110100001","1000000101001000","1000110100101011","1000101100011111","1000101011111111","0000000100000100","0000110100000110","1000011100010011","1001101000010001","1000110111011001","1000100001001001","1000011001101101","0000010010000000","1000010000011111","1000001000010111","1000101110111110","1000100011000110","0000010011100001","0000001001011101","0000110100111011","0000101000100011","0000100011101111","0000011001100100","0000001100011000","1001111101011010","1010010010000100","1000010110011000","0000010111110001","1000011001010100","1000010111110100","1000111111010101","1000110110110100","1000110001010100","1000000111100110","1000010111011110","1000010111001110","1000000111010000","1000100110000001","1000100101110100","1000000101011100","0000001100111000","1000010100010000","1000010100100111","1000000100110000","1000011100000100","0001000010101111","0000010000001100","0001000000111011","0000000000110100","1000111000010011","1001011101111100","1000010000001101","1000010000001010","1001000111010011","0000100100111000","1000001010011011","0000010010100101","0000000010001000","1000100000011111","1000001001101011","1000001100000100","1000001111010010","1000000010000100","1000010001110010","0000001111111101","0000011000001100","0000010010101001","0000010101001011","0000001101110011","0000000110101001","0000101111000110","1000101001100010","1000010101000101","0000010101011000","0000011010100011","0000110110010000","0000101010111110","0000001000000101","1000011111100010","0000010110011110","0000011011001001","0000011111100111","0000010010010101","0000000111010011","1000100000110100","1000000000010101","1000000001011001","1000101011001011","1000110010000101","1000001011001101","0000010101010101","0000011001111001","1000001111001011","1000001111000011","1000000001011100","0000001110100111","1000001010101100","0000100001001000","0000001100111011","1001000111110010","0000000101000000","1000011111111101","1000001000100110","1000000001101011","0000110000010011","0000110001010010","1000010100001101","1000010010110010","1000010110011111","0001010101110110","0000000110111011","0000001000101011","0000000101011101","0000001011000011","1000111111001010","1001010101011001","1001100110111000","1000101101100001","1000010011111011","1000010000000101","1000011100011100","1000000000000100","0000100000010100","0000100100111100","0001000000110011","0000010101110100","1001001000001001","1000100100000000","0000000001111011","0000010010001101","0001001001100011","1000000100111110","1000000010011100","0000000101100101","1001001000011010","1000100101100010","1000101101000001","0000110101011001","0000000000001001","1000010001010100","1000001000010101","1000001110101110","1000111101101111","1001000111110011","1000001000110010","1000010111011011","1001010110101100","1000010001010101","0000001101011110","0000010111010100","1000000011010111","1000100101010110","0000100001001101","1000011010110111","1000101011000101","1000101011110000","1000110010010110","1000000000011001","0001100101011010","0000000010000010","1000000000010111","0000000001101011","1000010001101001","1001001001101000","1001100001111001","1000011011000000","1000001010000011","1000011100000000","1000100111001011","1000011101010010","1000101111010101","1000111111011011","1000111110001101","1000111000011101","1001000101011110","1001000011111000","1001010111010001","1000011010000011","1000001011110111","1000010101111010","0000011110001101","1000000001011100","1000011100011101","1000100110111100","1001001000000101","0000001101101100","0000111000101000","0000000101011000","1000000010011111","1000000110100000","1000000101001110","1001000111101100","1010100000110100","1001010001000110","1001110111010000","1001010100011100","1000110001111000","1001100101100110","1011000101001010","1011001110111100","1001001111011010","1001101010111010","1001010110001110","1001111100011010","1100110000001111","1101000010000001","1110101110011111","1100001101100110","1011011011111101","1010000010101001","1001100001110111","1001001001110010","1000111101001110","1000010000111101","1000010000011110","0000000010000010","0000000010000100","0000000011100111","0000000001010110","1000100101001000","1001010100100101","1010001001011000","1001011001100011","1001100110100010","1011010010110010","1010011101011010","1010110001110110","1011000101101010","1011100011110000","1011011101100010","1010011111001111","1001011101000100","1010001101111101","1010110101011010","1010000000111000","1001101001011011","1010011100010101","1001101111010010","1001010110001100","1000110011000110","0000000001111011","1000000001101111","1000000110101001","1000000001011011","0000000001101010","0000000000111111","1000000100101110","0000000010001010","1000000000100010","1000001010111111","1000001011000011","1000000100110100","1000010110110010","1000011001110011","1000111100111101","1001101101101000","1001010111101010","1001101101100110","1001101011100001","1001000101111111","1000111101110110","1000111110100011","1000111010001100","1000110100100111","1000010010011001","1000011111110010","1000100110000111","1000010100001110","1000000001010111","0000000011011000","1000000010101110","1000000011001100");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
