library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity fully_connected_layer_0_3 is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_3 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end fully_connected_layer_0_3 ;
architecture Behavioral of fully_connected_layer_0_3 is
signal store_sum : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_0 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000100";
signal store_weight_0 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_1 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000110";
signal store_weight_1 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_2 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001000";
signal store_weight_2 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_3 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000010";
signal store_weight_3 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_4 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001100";
signal store_weight_4 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_5 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010101";
signal store_weight_5 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_6 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001100";
signal store_weight_6 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_7 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001011";
signal store_weight_7 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_8 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_8 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_9 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010101";
signal store_weight_9 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_10 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010100";
signal store_weight_10 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_11 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000001";
signal store_weight_11 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_12 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000100";
signal store_weight_12 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_13 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000001";
signal store_weight_13 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_14 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100111";
signal store_weight_14 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_15 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011100";
signal store_weight_15 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_16 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001111";
signal store_weight_16 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_17 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010101";
signal store_weight_17 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_18 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_18 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_19 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000000";
signal store_weight_19 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_20 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010110";
signal store_weight_20 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_21 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010011";
signal store_weight_21 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_22 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001000";
signal store_weight_22 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_23 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001111";
signal store_weight_23 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_24 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001010";
signal store_weight_24 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_25 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001000";
signal store_weight_25 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_26 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010010";
signal store_weight_26 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_27 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010010";
signal store_weight_27 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_28 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001011";
signal store_weight_28 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_29 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001111";
signal store_weight_29 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_30 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001101";
signal store_weight_30 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_31 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000010";
signal store_weight_31 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_32 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110101";
signal store_weight_32 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_33 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100100";
signal store_weight_33 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_34 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000111";
signal store_weight_34 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_35 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100001101";
signal store_weight_35 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_36 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100000101";
signal store_weight_36 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_37 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100100100";
signal store_weight_37 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_38 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101100110";
signal store_weight_38 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_39 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110111";
signal store_weight_39 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_40 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011100";
signal store_weight_40 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_41 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110110";
signal store_weight_41 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_42 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011011";
signal store_weight_42 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_43 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011010";
signal store_weight_43 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_44 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011001000";
signal store_weight_44 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_45 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100100";
signal store_weight_45 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_46 : STD_LOGIC_VECTOR(15 downto 0) := "1000001000101011";
signal store_weight_46 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_47 : STD_LOGIC_VECTOR(15 downto 0) := "1000001001100111";
signal store_weight_47 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_48 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110110011";
signal store_weight_48 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_49 : STD_LOGIC_VECTOR(15 downto 0) := "1000000111000111";
signal store_weight_49 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_50 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010111010";
signal store_weight_50 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_51 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010100011";
signal store_weight_51 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_52 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_52 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_53 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001100";
signal store_weight_53 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_54 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000101";
signal store_weight_54 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_55 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000110";
signal store_weight_55 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_56 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000001";
signal store_weight_56 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_57 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001101";
signal store_weight_57 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_58 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010010";
signal store_weight_58 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_59 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101001";
signal store_weight_59 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_60 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011000";
signal store_weight_60 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_61 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100001111";
signal store_weight_61 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_62 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011111";
signal store_weight_62 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_63 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011001";
signal store_weight_63 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_64 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010101101";
signal store_weight_64 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_65 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000011";
signal store_weight_65 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_66 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011100111";
signal store_weight_66 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_67 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011010000";
signal store_weight_67 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_68 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011010010";
signal store_weight_68 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_69 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100100";
signal store_weight_69 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_70 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000010";
signal store_weight_70 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_71 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011100001";
signal store_weight_71 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_72 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010101";
signal store_weight_72 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_73 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100111100";
signal store_weight_73 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_74 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100000101";
signal store_weight_74 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_75 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101000110";
signal store_weight_75 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_76 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010100010";
signal store_weight_76 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_77 : STD_LOGIC_VECTOR(15 downto 0) := "1000001001111101";
signal store_weight_77 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_78 : STD_LOGIC_VECTOR(15 downto 0) := "1000001000110000";
signal store_weight_78 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_79 : STD_LOGIC_VECTOR(15 downto 0) := "1000001000001000";
signal store_weight_79 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_80 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110000011";
signal store_weight_80 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_81 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001110";
signal store_weight_81 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_82 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001110";
signal store_weight_82 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_83 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001001";
signal store_weight_83 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_84 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010001";
signal store_weight_84 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_85 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_85 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_86 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001101";
signal store_weight_86 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_87 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011111";
signal store_weight_87 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_88 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100110";
signal store_weight_88 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_89 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011101100";
signal store_weight_89 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_90 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100110001";
signal store_weight_90 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_91 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100010111";
signal store_weight_91 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_92 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010101";
signal store_weight_92 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_93 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000110";
signal store_weight_93 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_94 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011101100";
signal store_weight_94 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_95 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101111110";
signal store_weight_95 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_96 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100001011";
signal store_weight_96 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_97 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100101001";
signal store_weight_97 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_98 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101001001";
signal store_weight_98 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_99 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101111100";
signal store_weight_99 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_100 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110010001";
signal store_weight_100 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_101 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110111011";
signal store_weight_101 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_102 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110101110";
signal store_weight_102 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_103 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101101000";
signal store_weight_103 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_104 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101010101";
signal store_weight_104 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_105 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010100011";
signal store_weight_105 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_106 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010110";
signal store_weight_106 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_107 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110011";
signal store_weight_107 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_108 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101000";
signal store_weight_108 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_109 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010100";
signal store_weight_109 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_110 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101001";
signal store_weight_110 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_111 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000101";
signal store_weight_111 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_112 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010000";
signal store_weight_112 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_113 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001011";
signal store_weight_113 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_114 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111011";
signal store_weight_114 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_115 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001010";
signal store_weight_115 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_116 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100100";
signal store_weight_116 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_117 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101000010";
signal store_weight_117 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_118 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011010000";
signal store_weight_118 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_119 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011001010";
signal store_weight_119 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_120 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101011";
signal store_weight_120 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_121 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100001";
signal store_weight_121 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_122 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011011";
signal store_weight_122 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_123 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100100";
signal store_weight_123 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_124 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111010";
signal store_weight_124 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_125 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101101";
signal store_weight_125 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_126 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000111";
signal store_weight_126 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_127 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000001";
signal store_weight_127 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_128 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111001";
signal store_weight_128 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_129 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000110";
signal store_weight_129 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_130 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101101";
signal store_weight_130 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_131 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110110";
signal store_weight_131 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_132 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111011";
signal store_weight_132 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_133 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011010100";
signal store_weight_133 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_134 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001110";
signal store_weight_134 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_135 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011001010";
signal store_weight_135 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_136 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011100";
signal store_weight_136 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_137 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010110";
signal store_weight_137 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_138 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101000";
signal store_weight_138 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_139 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110011";
signal store_weight_139 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_140 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001101";
signal store_weight_140 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_141 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001010";
signal store_weight_141 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_142 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101111";
signal store_weight_142 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_143 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011000111";
signal store_weight_143 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_144 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001011";
signal store_weight_144 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_145 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101111100";
signal store_weight_145 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_146 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010110110";
signal store_weight_146 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_147 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001000";
signal store_weight_147 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_148 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110011";
signal store_weight_148 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_149 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000111";
signal store_weight_149 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_150 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000101";
signal store_weight_150 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_151 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001011";
signal store_weight_151 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_152 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101101";
signal store_weight_152 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_153 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110010";
signal store_weight_153 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_154 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000101";
signal store_weight_154 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_155 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010001";
signal store_weight_155 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_156 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100010";
signal store_weight_156 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_157 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000111";
signal store_weight_157 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_158 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100101";
signal store_weight_158 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_159 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100100";
signal store_weight_159 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_160 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100100011";
signal store_weight_160 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_161 : STD_LOGIC_VECTOR(15 downto 0) := "0000000110001000";
signal store_weight_161 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_162 : STD_LOGIC_VECTOR(15 downto 0) := "0000000110011001";
signal store_weight_162 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_163 : STD_LOGIC_VECTOR(15 downto 0) := "0000000110110011";
signal store_weight_163 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_164 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101001100";
signal store_weight_164 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_165 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011101100";
signal store_weight_165 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_166 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011010010";
signal store_weight_166 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_167 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000000";
signal store_weight_167 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_168 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001111";
signal store_weight_168 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_169 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111110";
signal store_weight_169 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_170 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011110";
signal store_weight_170 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_171 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001011";
signal store_weight_171 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_172 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110100";
signal store_weight_172 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_173 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101011101";
signal store_weight_173 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_174 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011100011";
signal store_weight_174 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_175 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100011100";
signal store_weight_175 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_176 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100110001";
signal store_weight_176 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_177 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101010111";
signal store_weight_177 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_178 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100100011";
signal store_weight_178 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_179 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010000";
signal store_weight_179 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_180 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101011";
signal store_weight_180 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_181 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001000";
signal store_weight_181 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_182 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011001";
signal store_weight_182 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_183 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101000";
signal store_weight_183 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_184 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001011";
signal store_weight_184 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_185 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011111";
signal store_weight_185 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_186 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001101";
signal store_weight_186 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_187 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101110";
signal store_weight_187 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_188 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000001";
signal store_weight_188 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_189 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000111";
signal store_weight_189 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_190 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000010";
signal store_weight_190 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_191 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010100111";
signal store_weight_191 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_192 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101001";
signal store_weight_192 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_193 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100011101";
signal store_weight_193 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_194 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101001001";
signal store_weight_194 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_195 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011001111";
signal store_weight_195 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_196 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011100";
signal store_weight_196 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_197 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000101";
signal store_weight_197 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_198 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010000";
signal store_weight_198 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_199 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010011011";
signal store_weight_199 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_200 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101111101";
signal store_weight_200 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_201 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011011011";
signal store_weight_201 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_202 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100001100";
signal store_weight_202 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_203 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011111110";
signal store_weight_203 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_204 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100101100";
signal store_weight_204 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_205 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011100110";
signal store_weight_205 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_206 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000010";
signal store_weight_206 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_207 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010111";
signal store_weight_207 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_208 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_208 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_209 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111000";
signal store_weight_209 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_210 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110000";
signal store_weight_210 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_211 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100100";
signal store_weight_211 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_212 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000000";
signal store_weight_212 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_213 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001101";
signal store_weight_213 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_214 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010011";
signal store_weight_214 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_215 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010001";
signal store_weight_215 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_216 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101000";
signal store_weight_216 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_217 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000110";
signal store_weight_217 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_218 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000111";
signal store_weight_218 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_219 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100100";
signal store_weight_219 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_220 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110000";
signal store_weight_220 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_221 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101101";
signal store_weight_221 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_222 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110101";
signal store_weight_222 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_223 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011101110";
signal store_weight_223 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_224 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001101";
signal store_weight_224 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_225 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010100000";
signal store_weight_225 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_226 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111010";
signal store_weight_226 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_227 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011110000";
signal store_weight_227 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_228 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100111001";
signal store_weight_228 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_229 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010110111";
signal store_weight_229 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_230 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100011011";
signal store_weight_230 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_231 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100101";
signal store_weight_231 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_232 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101001";
signal store_weight_232 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_233 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000111";
signal store_weight_233 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_234 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110101";
signal store_weight_234 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_235 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001110";
signal store_weight_235 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_236 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011011";
signal store_weight_236 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_237 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101010";
signal store_weight_237 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_238 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000100";
signal store_weight_238 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_239 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001110";
signal store_weight_239 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_240 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101000";
signal store_weight_240 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_241 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010001";
signal store_weight_241 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_242 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111001";
signal store_weight_242 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_243 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011010";
signal store_weight_243 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_244 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111010";
signal store_weight_244 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_245 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010011";
signal store_weight_245 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_246 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110001";
signal store_weight_246 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_247 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101101";
signal store_weight_247 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_248 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001000";
signal store_weight_248 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_249 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111001";
signal store_weight_249 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_250 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010110";
signal store_weight_250 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_251 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100011110";
signal store_weight_251 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_252 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011001";
signal store_weight_252 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_253 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011001101";
signal store_weight_253 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_254 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000001";
signal store_weight_254 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_255 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011100010";
signal store_weight_255 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_256 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101011011";
signal store_weight_256 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_257 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011011001";
signal store_weight_257 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_258 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111011";
signal store_weight_258 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_259 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100101";
signal store_weight_259 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_260 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101011";
signal store_weight_260 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_261 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000101";
signal store_weight_261 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_262 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011000";
signal store_weight_262 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_263 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000111";
signal store_weight_263 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_264 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110000";
signal store_weight_264 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_265 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101100";
signal store_weight_265 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_266 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001101";
signal store_weight_266 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_267 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111001";
signal store_weight_267 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_268 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000111";
signal store_weight_268 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_269 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010011110";
signal store_weight_269 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_270 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001000";
signal store_weight_270 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_271 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110100";
signal store_weight_271 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_272 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110011";
signal store_weight_272 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_273 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000110";
signal store_weight_273 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_274 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_274 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_275 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010011";
signal store_weight_275 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_276 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001101";
signal store_weight_276 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_277 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110101";
signal store_weight_277 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_278 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011101011";
signal store_weight_278 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_279 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010101";
signal store_weight_279 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_280 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101000";
signal store_weight_280 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_281 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001001";
signal store_weight_281 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_282 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110000100";
signal store_weight_282 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_283 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100111100";
signal store_weight_283 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_284 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000111";
signal store_weight_284 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_285 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001101";
signal store_weight_285 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_286 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100111";
signal store_weight_286 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_287 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111111";
signal store_weight_287 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_288 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100111";
signal store_weight_288 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_289 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001101001";
signal store_weight_289 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_290 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000110";
signal store_weight_290 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_291 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111000";
signal store_weight_291 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_292 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011011100";
signal store_weight_292 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_293 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110010";
signal store_weight_293 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_294 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001001";
signal store_weight_294 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_295 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal store_weight_295 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_296 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010110000";
signal store_weight_296 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_297 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111011";
signal store_weight_297 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_298 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101001";
signal store_weight_298 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_299 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101110";
signal store_weight_299 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_300 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101001";
signal store_weight_300 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_301 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010100";
signal store_weight_301 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_302 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010011";
signal store_weight_302 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_303 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000101";
signal store_weight_303 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_304 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100011";
signal store_weight_304 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_305 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001000";
signal store_weight_305 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_306 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111110";
signal store_weight_306 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_307 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111111";
signal store_weight_307 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_308 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000000";
signal store_weight_308 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_309 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110100";
signal store_weight_309 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_310 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010111100";
signal store_weight_310 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_311 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100001000";
signal store_weight_311 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_312 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010101";
signal store_weight_312 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_313 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000011";
signal store_weight_313 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_314 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001100";
signal store_weight_314 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_315 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011000011";
signal store_weight_315 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_316 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111010";
signal store_weight_316 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_317 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111001";
signal store_weight_317 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_318 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111110";
signal store_weight_318 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_319 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111011";
signal store_weight_319 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_320 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100010";
signal store_weight_320 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_321 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000011";
signal store_weight_321 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_322 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110110";
signal store_weight_322 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_323 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000100";
signal store_weight_323 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_324 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000110";
signal store_weight_324 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_325 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011011011";
signal store_weight_325 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_326 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000110";
signal store_weight_326 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_327 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101111";
signal store_weight_327 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_328 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011001";
signal store_weight_328 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_329 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010000";
signal store_weight_329 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_330 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010000";
signal store_weight_330 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_331 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100111";
signal store_weight_331 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_332 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000101";
signal store_weight_332 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_333 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101010";
signal store_weight_333 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_334 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011011001";
signal store_weight_334 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_335 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001001";
signal store_weight_335 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_336 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000101";
signal store_weight_336 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_337 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011110010";
signal store_weight_337 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_338 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011001011";
signal store_weight_338 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_339 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100110";
signal store_weight_339 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_340 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010011110";
signal store_weight_340 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_341 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100111";
signal store_weight_341 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_342 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100110";
signal store_weight_342 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_343 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010011";
signal store_weight_343 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_344 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110100";
signal store_weight_344 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_345 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101111";
signal store_weight_345 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_346 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111000";
signal store_weight_346 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_347 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010101";
signal store_weight_347 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_348 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010100101";
signal store_weight_348 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_349 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100110001";
signal store_weight_349 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_350 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011110111";
signal store_weight_350 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_351 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110100";
signal store_weight_351 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_352 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011110100";
signal store_weight_352 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_353 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010011100";
signal store_weight_353 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_354 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010011";
signal store_weight_354 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_355 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011110";
signal store_weight_355 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_356 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101101";
signal store_weight_356 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_357 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100011";
signal store_weight_357 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_358 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001111";
signal store_weight_358 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_359 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100100";
signal store_weight_359 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_360 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100001";
signal store_weight_360 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_361 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010000";
signal store_weight_361 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_362 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011010010";
signal store_weight_362 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_363 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110000";
signal store_weight_363 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_364 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010100";
signal store_weight_364 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_365 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100000";
signal store_weight_365 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_366 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011010111";
signal store_weight_366 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_367 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111100";
signal store_weight_367 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_368 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101100";
signal store_weight_368 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_369 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010110";
signal store_weight_369 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_370 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010111";
signal store_weight_370 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_371 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_371 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_372 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_372 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_373 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000101";
signal store_weight_373 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_374 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010110";
signal store_weight_374 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_375 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011000110";
signal store_weight_375 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_376 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011111010";
signal store_weight_376 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_377 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101010110";
signal store_weight_377 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_378 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011100111";
signal store_weight_378 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_379 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000110";
signal store_weight_379 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_380 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010101011";
signal store_weight_380 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_381 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110110";
signal store_weight_381 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_382 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111000";
signal store_weight_382 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_383 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111110";
signal store_weight_383 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_384 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011001";
signal store_weight_384 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_385 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000010";
signal store_weight_385 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_386 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011011";
signal store_weight_386 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_387 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001111";
signal store_weight_387 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_388 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100010";
signal store_weight_388 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_389 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001001";
signal store_weight_389 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_390 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100111010";
signal store_weight_390 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_391 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101101";
signal store_weight_391 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_392 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010110";
signal store_weight_392 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_393 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100101100";
signal store_weight_393 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_394 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011011101";
signal store_weight_394 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_395 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010011001";
signal store_weight_395 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_396 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010001";
signal store_weight_396 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_397 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000101";
signal store_weight_397 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_398 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001011";
signal store_weight_398 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_399 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000011";
signal store_weight_399 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_400 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010100";
signal store_weight_400 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_401 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011110";
signal store_weight_401 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_402 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001101111";
signal store_weight_402 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_403 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111100";
signal store_weight_403 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_404 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101010010";
signal store_weight_404 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_405 : STD_LOGIC_VECTOR(15 downto 0) := "0000000110101000";
signal store_weight_405 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_406 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011100010";
signal store_weight_406 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_407 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110000";
signal store_weight_407 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_408 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001000";
signal store_weight_408 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_409 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011001101";
signal store_weight_409 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_410 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010100";
signal store_weight_410 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_411 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101110";
signal store_weight_411 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_412 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111010";
signal store_weight_412 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_413 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010001";
signal store_weight_413 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_414 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000111";
signal store_weight_414 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_415 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110001";
signal store_weight_415 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_416 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101101";
signal store_weight_416 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_417 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001100";
signal store_weight_417 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_418 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101010010";
signal store_weight_418 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_419 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011011101";
signal store_weight_419 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_420 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011101";
signal store_weight_420 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_421 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111111";
signal store_weight_421 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_422 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011101";
signal store_weight_422 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_423 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010101001";
signal store_weight_423 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_424 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100001";
signal store_weight_424 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_425 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001010";
signal store_weight_425 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_426 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111000";
signal store_weight_426 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_427 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101001";
signal store_weight_427 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_428 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011100";
signal store_weight_428 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_429 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101111";
signal store_weight_429 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_430 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001010111";
signal store_weight_430 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_431 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111010";
signal store_weight_431 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_432 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011011111";
signal store_weight_432 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_433 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011110101";
signal store_weight_433 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_434 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110100";
signal store_weight_434 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_435 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000001";
signal store_weight_435 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_436 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001000";
signal store_weight_436 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_437 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000111";
signal store_weight_437 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_438 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010111000";
signal store_weight_438 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_439 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000100";
signal store_weight_439 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_440 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010011101";
signal store_weight_440 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_441 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000100";
signal store_weight_441 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_442 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000011";
signal store_weight_442 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_443 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111100";
signal store_weight_443 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_444 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101010";
signal store_weight_444 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_445 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000110";
signal store_weight_445 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_446 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011001010";
signal store_weight_446 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_447 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101100";
signal store_weight_447 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_448 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001000";
signal store_weight_448 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_449 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010111100";
signal store_weight_449 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_450 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011011";
signal store_weight_450 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_451 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111111";
signal store_weight_451 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_452 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000100";
signal store_weight_452 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_453 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100111";
signal store_weight_453 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_454 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110000";
signal store_weight_454 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_455 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010000";
signal store_weight_455 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_456 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010001";
signal store_weight_456 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_457 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000011";
signal store_weight_457 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_458 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111101";
signal store_weight_458 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_459 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110011";
signal store_weight_459 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_460 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010110001";
signal store_weight_460 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_461 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100110";
signal store_weight_461 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_462 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110000";
signal store_weight_462 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_463 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000110";
signal store_weight_463 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_464 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100011";
signal store_weight_464 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_465 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100101";
signal store_weight_465 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_466 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001000";
signal store_weight_466 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_467 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110111";
signal store_weight_467 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_468 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001111";
signal store_weight_468 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_469 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101000";
signal store_weight_469 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_470 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111100";
signal store_weight_470 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_471 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000100";
signal store_weight_471 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_472 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001101";
signal store_weight_472 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_473 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010111";
signal store_weight_473 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_474 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011001100";
signal store_weight_474 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_475 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100100000";
signal store_weight_475 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_476 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001011";
signal store_weight_476 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_477 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010101";
signal store_weight_477 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_478 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001101";
signal store_weight_478 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_479 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010101111";
signal store_weight_479 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_480 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001101";
signal store_weight_480 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_481 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110000";
signal store_weight_481 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_482 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001010010";
signal store_weight_482 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_483 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010110";
signal store_weight_483 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_484 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011101";
signal store_weight_484 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_485 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001010";
signal store_weight_485 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_486 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001100";
signal store_weight_486 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_487 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111000";
signal store_weight_487 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_488 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000010";
signal store_weight_488 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_489 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000100";
signal store_weight_489 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_490 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001100";
signal store_weight_490 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_491 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011111";
signal store_weight_491 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_492 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011010";
signal store_weight_492 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_493 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100011";
signal store_weight_493 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_494 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010101010";
signal store_weight_494 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_495 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010011";
signal store_weight_495 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_496 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111100";
signal store_weight_496 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_497 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110011";
signal store_weight_497 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_498 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101011";
signal store_weight_498 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_499 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111010";
signal store_weight_499 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_500 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011001";
signal store_weight_500 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_501 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000100";
signal store_weight_501 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_502 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001111";
signal store_weight_502 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_503 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011100000";
signal store_weight_503 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_504 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011010";
signal store_weight_504 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_505 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011011000";
signal store_weight_505 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_506 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100000010";
signal store_weight_506 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_507 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110011";
signal store_weight_507 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_508 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111000";
signal store_weight_508 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_509 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010110101";
signal store_weight_509 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_510 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001100";
signal store_weight_510 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_511 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011110";
signal store_weight_511 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_512 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111000";
signal store_weight_512 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_513 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111000";
signal store_weight_513 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_514 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010010";
signal store_weight_514 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_515 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011111";
signal store_weight_515 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_516 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001010";
signal store_weight_516 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_517 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011110";
signal store_weight_517 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_518 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000100";
signal store_weight_518 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_519 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001101110";
signal store_weight_519 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_520 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110110";
signal store_weight_520 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_521 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001100";
signal store_weight_521 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_522 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001011";
signal store_weight_522 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_523 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100011";
signal store_weight_523 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_524 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000011";
signal store_weight_524 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_525 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100011";
signal store_weight_525 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_526 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010101";
signal store_weight_526 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_527 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000101";
signal store_weight_527 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_528 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110100";
signal store_weight_528 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_529 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111111";
signal store_weight_529 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_530 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110100";
signal store_weight_530 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_531 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011110001";
signal store_weight_531 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_532 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000101";
signal store_weight_532 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_533 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000110";
signal store_weight_533 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_534 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011010111";
signal store_weight_534 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_535 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100111";
signal store_weight_535 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_536 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110000";
signal store_weight_536 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_537 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001110";
signal store_weight_537 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_538 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010101";
signal store_weight_538 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_539 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100100";
signal store_weight_539 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_540 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011010111";
signal store_weight_540 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_541 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001101010";
signal store_weight_541 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_542 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100011";
signal store_weight_542 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_543 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100000";
signal store_weight_543 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_544 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110001";
signal store_weight_544 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_545 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101010";
signal store_weight_545 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_546 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000101";
signal store_weight_546 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_547 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011010";
signal store_weight_547 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_548 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111101";
signal store_weight_548 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_549 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010001";
signal store_weight_549 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_550 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010101";
signal store_weight_550 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_551 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110101";
signal store_weight_551 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_552 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011110";
signal store_weight_552 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_553 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000111";
signal store_weight_553 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_554 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001011";
signal store_weight_554 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_555 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100101001";
signal store_weight_555 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_556 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111110";
signal store_weight_556 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_557 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111100";
signal store_weight_557 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_558 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101010011";
signal store_weight_558 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_559 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111101";
signal store_weight_559 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_560 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000001";
signal store_weight_560 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_561 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001111";
signal store_weight_561 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_562 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001101";
signal store_weight_562 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_563 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100010110";
signal store_weight_563 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_564 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_564 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_565 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011101";
signal store_weight_565 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_566 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100000";
signal store_weight_566 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_567 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001001";
signal store_weight_567 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_568 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010111";
signal store_weight_568 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_569 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111100";
signal store_weight_569 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_570 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001010";
signal store_weight_570 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_571 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010010";
signal store_weight_571 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_572 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111101";
signal store_weight_572 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_573 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010001";
signal store_weight_573 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_574 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010110001";
signal store_weight_574 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_575 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010111";
signal store_weight_575 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_576 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011100";
signal store_weight_576 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_577 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100010";
signal store_weight_577 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_578 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101000";
signal store_weight_578 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_579 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011100";
signal store_weight_579 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_580 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100111";
signal store_weight_580 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_581 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111111";
signal store_weight_581 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_582 : STD_LOGIC_VECTOR(15 downto 0) := "0000000110000010";
signal store_weight_582 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_583 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101011";
signal store_weight_583 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_584 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011110011";
signal store_weight_584 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_585 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000011";
signal store_weight_585 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_586 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111011";
signal store_weight_586 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_587 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001101000";
signal store_weight_587 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_588 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010001";
signal store_weight_588 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_589 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111000";
signal store_weight_589 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_590 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010101001";
signal store_weight_590 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_591 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111100";
signal store_weight_591 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_592 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110011";
signal store_weight_592 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_593 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100110";
signal store_weight_593 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_594 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000111010";
signal store_weight_594 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_595 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001001";
signal store_weight_595 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_596 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011011";
signal store_weight_596 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_597 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001011";
signal store_weight_597 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_598 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111001";
signal store_weight_598 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_599 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010010";
signal store_weight_599 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_600 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100011";
signal store_weight_600 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_601 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111100";
signal store_weight_601 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_602 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010110";
signal store_weight_602 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_603 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100001";
signal store_weight_603 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_604 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010111";
signal store_weight_604 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_605 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101111";
signal store_weight_605 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_606 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101101";
signal store_weight_606 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_607 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011101";
signal store_weight_607 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_608 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011010000";
signal store_weight_608 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_609 : STD_LOGIC_VECTOR(15 downto 0) := "0000000111100100";
signal store_weight_609 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_610 : STD_LOGIC_VECTOR(15 downto 0) := "0000001000010110";
signal store_weight_610 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_611 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101110011";
signal store_weight_611 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_612 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111011";
signal store_weight_612 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_613 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101010";
signal store_weight_613 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_614 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100011";
signal store_weight_614 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_615 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001100";
signal store_weight_615 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_616 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110010";
signal store_weight_616 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_617 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011011";
signal store_weight_617 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_618 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011001011";
signal store_weight_618 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_619 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011000";
signal store_weight_619 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_620 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100100";
signal store_weight_620 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_621 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011110";
signal store_weight_621 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_622 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111111";
signal store_weight_622 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_623 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101000";
signal store_weight_623 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_624 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000001";
signal store_weight_624 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_625 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001000";
signal store_weight_625 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_626 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111000";
signal store_weight_626 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_627 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110000";
signal store_weight_627 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_628 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010000";
signal store_weight_628 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_629 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000101000";
signal store_weight_629 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_630 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000000";
signal store_weight_630 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_631 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100000";
signal store_weight_631 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_632 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011101";
signal store_weight_632 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_633 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001011";
signal store_weight_633 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_634 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111100";
signal store_weight_634 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_635 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111001";
signal store_weight_635 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_636 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011110000";
signal store_weight_636 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_637 : STD_LOGIC_VECTOR(15 downto 0) := "0000000110110011";
signal store_weight_637 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_638 : STD_LOGIC_VECTOR(15 downto 0) := "0000000110010110";
signal store_weight_638 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_639 : STD_LOGIC_VECTOR(15 downto 0) := "0000001000110010";
signal store_weight_639 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_640 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100110110";
signal store_weight_640 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_641 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011101000";
signal store_weight_641 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_642 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110111";
signal store_weight_642 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_643 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001011";
signal store_weight_643 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_644 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001010";
signal store_weight_644 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_645 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000101";
signal store_weight_645 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_646 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000111";
signal store_weight_646 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_647 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010000";
signal store_weight_647 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_648 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011010110";
signal store_weight_648 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_649 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101011";
signal store_weight_649 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_650 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100000100";
signal store_weight_650 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_651 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010101";
signal store_weight_651 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_652 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010001";
signal store_weight_652 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_653 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001000";
signal store_weight_653 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_654 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110011";
signal store_weight_654 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_655 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000110100";
signal store_weight_655 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_656 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111010";
signal store_weight_656 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_657 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010100011";
signal store_weight_657 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_658 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011101";
signal store_weight_658 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_659 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010010100";
signal store_weight_659 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_660 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111011";
signal store_weight_660 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_661 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001011101";
signal store_weight_661 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_662 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000110";
signal store_weight_662 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_663 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100100";
signal store_weight_663 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_664 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011010100";
signal store_weight_664 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_665 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011000101";
signal store_weight_665 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_666 : STD_LOGIC_VECTOR(15 downto 0) := "0000000100100010";
signal store_weight_666 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_667 : STD_LOGIC_VECTOR(15 downto 0) := "0000000101111100";
signal store_weight_667 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_668 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101110";
signal store_weight_668 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_669 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101001";
signal store_weight_669 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_670 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000110";
signal store_weight_670 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_671 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000010";
signal store_weight_671 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_672 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000111";
signal store_weight_672 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_673 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000001";
signal store_weight_673 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_674 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100100";
signal store_weight_674 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_675 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011100";
signal store_weight_675 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_676 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101010";
signal store_weight_676 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_677 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011110110";
signal store_weight_677 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_678 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011010011";
signal store_weight_678 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_679 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010010111";
signal store_weight_679 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_680 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001101";
signal store_weight_680 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_681 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101000";
signal store_weight_681 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_682 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100011";
signal store_weight_682 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_683 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011011";
signal store_weight_683 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_684 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011110";
signal store_weight_684 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_685 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001011";
signal store_weight_685 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_686 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000100";
signal store_weight_686 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_687 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110000";
signal store_weight_687 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_688 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001110";
signal store_weight_688 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_689 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100101";
signal store_weight_689 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_690 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001100110";
signal store_weight_690 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_691 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010100110";
signal store_weight_691 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_692 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001111";
signal store_weight_692 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_693 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011100111";
signal store_weight_693 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_694 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010111011";
signal store_weight_694 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_695 : STD_LOGIC_VECTOR(15 downto 0) := "0000000111001111";
signal store_weight_695 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_696 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011111100";
signal store_weight_696 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_697 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001011";
signal store_weight_697 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_698 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000010";
signal store_weight_698 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_699 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001100";
signal store_weight_699 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_700 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001111";
signal store_weight_700 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_701 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000101";
signal store_weight_701 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_702 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010001101";
signal store_weight_702 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_703 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100001";
signal store_weight_703 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_704 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001000";
signal store_weight_704 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_705 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001110";
signal store_weight_705 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_706 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001011";
signal store_weight_706 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_707 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000110100";
signal store_weight_707 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_708 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000010";
signal store_weight_708 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_709 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal store_weight_709 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_710 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010101001";
signal store_weight_710 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_711 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000111";
signal store_weight_711 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_712 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100010";
signal store_weight_712 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_713 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111010";
signal store_weight_713 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_714 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001111010";
signal store_weight_714 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_715 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011011";
signal store_weight_715 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_716 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010001";
signal store_weight_716 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_717 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001111";
signal store_weight_717 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_718 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000100000";
signal store_weight_718 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_719 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001100";
signal store_weight_719 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_720 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000101";
signal store_weight_720 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_721 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011001011";
signal store_weight_721 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_722 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011110";
signal store_weight_722 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_723 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000000";
signal store_weight_723 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_724 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011001";
signal store_weight_724 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_725 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010011111";
signal store_weight_725 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_726 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001011";
signal store_weight_726 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_727 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010001";
signal store_weight_727 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_728 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001010";
signal store_weight_728 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_729 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010101";
signal store_weight_729 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_730 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000101";
signal store_weight_730 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_731 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001101000";
signal store_weight_731 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_732 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010100111";
signal store_weight_732 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_733 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011111";
signal store_weight_733 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_734 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010101";
signal store_weight_734 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_735 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000010";
signal store_weight_735 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_736 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000011111";
signal store_weight_736 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_737 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001110001";
signal store_weight_737 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_738 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010110";
signal store_weight_738 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_739 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001101000";
signal store_weight_739 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_740 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011001010";
signal store_weight_740 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_741 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000001";
signal store_weight_741 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_742 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001001000";
signal store_weight_742 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_743 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000111111";
signal store_weight_743 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_744 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000000";
signal store_weight_744 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_745 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000111";
signal store_weight_745 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_746 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001100001";
signal store_weight_746 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_747 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011001";
signal store_weight_747 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_748 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001111";
signal store_weight_748 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_749 : STD_LOGIC_VECTOR(15 downto 0) := "0000000001000001";
signal store_weight_749 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_750 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010111";
signal store_weight_750 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_751 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011011100";
signal store_weight_751 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_752 : STD_LOGIC_VECTOR(15 downto 0) := "0000000010000101";
signal store_weight_752 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_753 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001011000";
signal store_weight_753 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_754 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000010011";
signal store_weight_754 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_755 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000110";
signal store_weight_755 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_756 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000011";
signal store_weight_756 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_757 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001001";
signal store_weight_757 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_758 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010010";
signal store_weight_758 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_759 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000110";
signal store_weight_759 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_760 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010101110";
signal store_weight_760 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_761 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011111010";
signal store_weight_761 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_762 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000100000";
signal store_weight_762 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_763 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001111";
signal store_weight_763 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_764 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001001110";
signal store_weight_764 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_765 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000101000";
signal store_weight_765 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_766 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001010101";
signal store_weight_766 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_767 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000011100";
signal store_weight_767 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_768 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101110";
signal store_weight_768 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_769 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110101110";
signal store_weight_769 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_770 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001110001";
signal store_weight_770 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_771 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001110";
signal store_weight_771 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_772 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100010010";
signal store_weight_772 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_773 : STD_LOGIC_VECTOR(15 downto 0) := "1000000110000010";
signal store_weight_773 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_774 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010001101";
signal store_weight_774 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_775 : STD_LOGIC_VECTOR(15 downto 0) := "1000000010000011";
signal store_weight_775 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_776 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001000101";
signal store_weight_776 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_777 : STD_LOGIC_VECTOR(15 downto 0) := "1000000001101000";
signal store_weight_777 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_778 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010010";
signal store_weight_778 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_779 : STD_LOGIC_VECTOR(15 downto 0) := "1000000011000010";
signal store_weight_779 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_780 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000001110";
signal store_weight_780 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_781 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000011";
signal store_weight_781 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_782 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000001000";
signal store_weight_782 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_783 : STD_LOGIC_VECTOR(15 downto 0) := "1000000000010010";
signal store_weight_783 : STD_LOGIC_VECTOR(15 downto 0) ;
signal sum_0 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_1 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_2 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_3 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_4 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_5 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_6 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_7 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_8 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_9 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_10 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_11 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_12 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_13 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_14 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_15 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_16 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_17 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_18 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_19 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_20 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_21 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_22 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_23 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_24 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_25 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_26 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_27 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_28 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_29 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_30 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_31 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_32 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_33 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_34 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_35 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_36 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_37 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_38 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_39 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_40 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_41 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_42 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_43 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_44 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_45 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_46 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_47 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_48 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_49 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_50 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_51 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_52 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_53 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_54 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_55 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_56 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_57 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_58 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_59 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_60 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_61 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_62 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_63 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_64 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_65 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_66 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_67 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_68 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_69 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_70 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_71 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_72 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_73 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_74 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_75 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_76 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_77 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_78 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_79 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_80 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_81 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_82 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_83 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_84 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_85 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_86 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_87 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_88 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_89 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_90 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_91 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_92 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_93 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_94 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_95 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_96 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_97 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_98 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_99 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_100 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_101 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_102 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_103 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_104 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_105 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_106 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_107 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_108 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_109 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_110 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_111 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_112 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_113 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_114 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_115 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_116 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_117 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_118 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_119 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_120 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_121 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_122 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_123 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_124 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_125 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_126 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_127 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_128 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_129 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_130 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_131 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_132 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_133 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_134 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_135 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_136 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_137 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_138 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_139 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_140 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_141 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_142 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_143 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_144 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_145 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_146 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_147 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_148 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_149 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_150 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_151 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_152 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_153 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_154 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_155 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_156 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_157 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_158 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_159 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_160 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_161 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_162 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_163 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_164 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_165 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_166 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_167 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_168 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_169 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_170 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_171 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_172 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_173 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_174 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_175 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_176 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_177 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_178 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_179 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_180 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_181 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_182 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_183 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_184 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_185 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_186 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_187 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_188 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_189 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_190 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_191 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_192 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_193 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_194 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_195 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_196 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_197 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_198 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_199 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_200 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_201 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_202 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_203 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_204 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_205 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_206 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_207 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_208 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_209 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_210 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_211 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_212 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_213 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_214 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_215 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_216 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_217 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_218 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_219 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_220 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_221 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_222 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_223 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_224 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_225 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_226 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_227 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_228 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_229 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_230 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_231 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_232 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_233 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_234 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_235 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_236 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_237 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_238 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_239 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_240 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_241 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_242 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_243 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_244 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_245 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_246 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_247 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_248 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_249 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_250 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_251 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_252 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_253 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_254 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_255 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_256 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_257 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_258 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_259 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_260 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_261 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_262 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_263 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_264 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_265 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_266 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_267 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_268 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_269 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_270 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_271 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_272 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_273 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_274 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_275 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_276 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_277 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_278 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_279 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_280 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_281 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_282 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_283 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_284 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_285 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_286 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_287 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_288 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_289 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_290 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_291 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_292 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_293 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_294 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_295 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_296 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_297 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_298 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_299 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_300 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_301 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_302 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_303 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_304 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_305 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_306 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_307 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_308 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_309 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_310 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_311 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_312 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_313 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_314 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_315 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_316 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_317 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_318 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_319 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_320 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_321 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_322 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_323 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_324 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_325 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_326 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_327 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_328 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_329 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_330 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_331 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_332 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_333 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_334 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_335 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_336 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_337 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_338 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_339 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_340 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_341 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_342 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_343 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_344 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_345 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_346 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_347 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_348 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_349 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_350 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_351 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_352 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_353 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_354 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_355 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_356 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_357 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_358 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_359 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_360 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_361 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_362 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_363 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_364 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_365 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_366 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_367 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_368 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_369 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_370 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_371 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_372 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_373 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_374 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_375 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_376 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_377 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_378 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_379 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_380 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_381 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_382 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_383 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_384 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_385 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_386 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_387 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_388 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_389 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_390 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_391 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_392 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_393 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_394 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_395 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_396 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_397 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_398 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_399 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_400 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_401 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_402 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_403 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_404 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_405 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_406 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_407 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_408 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_409 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_410 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_411 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_412 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_413 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_414 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_415 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_416 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_417 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_418 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_419 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_420 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_421 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_422 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_423 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_424 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_425 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_426 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_427 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_428 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_429 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_430 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_431 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_432 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_433 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_434 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_435 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_436 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_437 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_438 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_439 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_440 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_441 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_442 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_443 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_444 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_445 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_446 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_447 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_448 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_449 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_450 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_451 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_452 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_453 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_454 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_455 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_456 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_457 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_458 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_459 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_460 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_461 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_462 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_463 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_464 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_465 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_466 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_467 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_468 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_469 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_470 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_471 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_472 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_473 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_474 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_475 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_476 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_477 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_478 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_479 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_480 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_481 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_482 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_483 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_484 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_485 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_486 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_487 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_488 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_489 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_490 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_491 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_492 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_493 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_494 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_495 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_496 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_497 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_498 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_499 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_500 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_501 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_502 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_503 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_504 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_505 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_506 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_507 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_508 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_509 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_510 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_511 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_512 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_513 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_514 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_515 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_516 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_517 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_518 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_519 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_520 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_521 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_522 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_523 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_524 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_525 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_526 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_527 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_528 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_529 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_530 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_531 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_532 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_533 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_534 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_535 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_536 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_537 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_538 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_539 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_540 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_541 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_542 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_543 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_544 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_545 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_546 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_547 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_548 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_549 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_550 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_551 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_552 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_553 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_554 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_555 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_556 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_557 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_558 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_559 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_560 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_561 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_562 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_563 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_564 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_565 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_566 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_567 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_568 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_569 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_570 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_571 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_572 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_573 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_574 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_575 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_576 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_577 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_578 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_579 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_580 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_581 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_582 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_583 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_584 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_585 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_586 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_587 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_588 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_589 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_590 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_591 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_592 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_593 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_594 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_595 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_596 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_597 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_598 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_599 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_600 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_601 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_602 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_603 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_604 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_605 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_606 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_607 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_608 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_609 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_610 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_611 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_612 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_613 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_614 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_615 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_616 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_617 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_618 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_619 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_620 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_621 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_622 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_623 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_624 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_625 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_626 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_627 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_628 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_629 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_630 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_631 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_632 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_633 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_634 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_635 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_636 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_637 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_638 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_639 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_640 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_641 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_642 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_643 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_644 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_645 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_646 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_647 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_648 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_649 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_650 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_651 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_652 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_653 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_654 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_655 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_656 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_657 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_658 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_659 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_660 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_661 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_662 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_663 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_664 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_665 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_666 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_667 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_668 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_669 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_670 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_671 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_672 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_673 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_674 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_675 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_676 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_677 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_678 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_679 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_680 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_681 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_682 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_683 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_684 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_685 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_686 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_687 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_688 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_689 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_690 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_691 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_692 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_693 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_694 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_695 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_696 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_697 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_698 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_699 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_700 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_701 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_702 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_703 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_704 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_705 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_706 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_707 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_708 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_709 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_710 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_711 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_712 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_713 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_714 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_715 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_716 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_717 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_718 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_719 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_720 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_721 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_722 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_723 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_724 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_725 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_726 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_727 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_728 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_729 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_730 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_731 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_732 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_733 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_734 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_735 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_736 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_737 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_738 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_739 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_740 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_741 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_742 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_743 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_744 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_745 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_746 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_747 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_748 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_749 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_750 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_751 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_752 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_753 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_754 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_755 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_756 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_757 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_758 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_759 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_760 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_761 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_762 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_763 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_764 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_765 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_766 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_767 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_768 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_769 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_770 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_771 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_772 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_773 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_774 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_775 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_776 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_777 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_778 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_779 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_780 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_781 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_782 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal biases : STD_LOGIC_VECTOR(15 downto 0) := "1000000000000011";
component  sigmoid is
	port (
		num:in integer ;
		y: out STD_LOGIC_VECTOR(15 downto 0)
		);
end component sigmoid;

component  nn_addition is
	Port (
		inputx : in STD_LOGIC_VECTOR(15 downto 0);
		inputy : in STD_LOGIC_VECTOR(15 downto 0);
		output : out STD_LOGIC_VECTOR(15 downto 0));
end component nn_addition;

component  nn_multiplication is
	Port (
		inputx : in STD_LOGIC_VECTOR(15 downto 0);
		inputy : in STD_LOGIC_VECTOR(15 downto 0);
		output : out STD_LOGIC_VECTOR(15 downto 0));
end component nn_multiplication;
begin
ut0_nn_multiplication: nn_multiplication port map(weight_0 , x_0 ,store_weight_0 );
ut1_nn_multiplication: nn_multiplication port map(weight_1 , x_1 ,store_weight_1 );
ut2_nn_multiplication: nn_multiplication port map(weight_2 , x_2 ,store_weight_2 );
ut3_nn_multiplication: nn_multiplication port map(weight_3 , x_3 ,store_weight_3 );
ut4_nn_multiplication: nn_multiplication port map(weight_4 , x_4 ,store_weight_4 );
ut5_nn_multiplication: nn_multiplication port map(weight_5 , x_5 ,store_weight_5 );
ut6_nn_multiplication: nn_multiplication port map(weight_6 , x_6 ,store_weight_6 );
ut7_nn_multiplication: nn_multiplication port map(weight_7 , x_7 ,store_weight_7 );
ut8_nn_multiplication: nn_multiplication port map(weight_8 , x_8 ,store_weight_8 );
ut9_nn_multiplication: nn_multiplication port map(weight_9 , x_9 ,store_weight_9 );
ut10_nn_multiplication: nn_multiplication port map(weight_10 , x_10 ,store_weight_10 );
ut11_nn_multiplication: nn_multiplication port map(weight_11 , x_11 ,store_weight_11 );
ut12_nn_multiplication: nn_multiplication port map(weight_12 , x_12 ,store_weight_12 );
ut13_nn_multiplication: nn_multiplication port map(weight_13 , x_13 ,store_weight_13 );
ut14_nn_multiplication: nn_multiplication port map(weight_14 , x_14 ,store_weight_14 );
ut15_nn_multiplication: nn_multiplication port map(weight_15 , x_15 ,store_weight_15 );
ut16_nn_multiplication: nn_multiplication port map(weight_16 , x_16 ,store_weight_16 );
ut17_nn_multiplication: nn_multiplication port map(weight_17 , x_17 ,store_weight_17 );
ut18_nn_multiplication: nn_multiplication port map(weight_18 , x_18 ,store_weight_18 );
ut19_nn_multiplication: nn_multiplication port map(weight_19 , x_19 ,store_weight_19 );
ut20_nn_multiplication: nn_multiplication port map(weight_20 , x_20 ,store_weight_20 );
ut21_nn_multiplication: nn_multiplication port map(weight_21 , x_21 ,store_weight_21 );
ut22_nn_multiplication: nn_multiplication port map(weight_22 , x_22 ,store_weight_22 );
ut23_nn_multiplication: nn_multiplication port map(weight_23 , x_23 ,store_weight_23 );
ut24_nn_multiplication: nn_multiplication port map(weight_24 , x_24 ,store_weight_24 );
ut25_nn_multiplication: nn_multiplication port map(weight_25 , x_25 ,store_weight_25 );
ut26_nn_multiplication: nn_multiplication port map(weight_26 , x_26 ,store_weight_26 );
ut27_nn_multiplication: nn_multiplication port map(weight_27 , x_27 ,store_weight_27 );
ut28_nn_multiplication: nn_multiplication port map(weight_28 , x_28 ,store_weight_28 );
ut29_nn_multiplication: nn_multiplication port map(weight_29 , x_29 ,store_weight_29 );
ut30_nn_multiplication: nn_multiplication port map(weight_30 , x_30 ,store_weight_30 );
ut31_nn_multiplication: nn_multiplication port map(weight_31 , x_31 ,store_weight_31 );
ut32_nn_multiplication: nn_multiplication port map(weight_32 , x_32 ,store_weight_32 );
ut33_nn_multiplication: nn_multiplication port map(weight_33 , x_33 ,store_weight_33 );
ut34_nn_multiplication: nn_multiplication port map(weight_34 , x_34 ,store_weight_34 );
ut35_nn_multiplication: nn_multiplication port map(weight_35 , x_35 ,store_weight_35 );
ut36_nn_multiplication: nn_multiplication port map(weight_36 , x_36 ,store_weight_36 );
ut37_nn_multiplication: nn_multiplication port map(weight_37 , x_37 ,store_weight_37 );
ut38_nn_multiplication: nn_multiplication port map(weight_38 , x_38 ,store_weight_38 );
ut39_nn_multiplication: nn_multiplication port map(weight_39 , x_39 ,store_weight_39 );
ut40_nn_multiplication: nn_multiplication port map(weight_40 , x_40 ,store_weight_40 );
ut41_nn_multiplication: nn_multiplication port map(weight_41 , x_41 ,store_weight_41 );
ut42_nn_multiplication: nn_multiplication port map(weight_42 , x_42 ,store_weight_42 );
ut43_nn_multiplication: nn_multiplication port map(weight_43 , x_43 ,store_weight_43 );
ut44_nn_multiplication: nn_multiplication port map(weight_44 , x_44 ,store_weight_44 );
ut45_nn_multiplication: nn_multiplication port map(weight_45 , x_45 ,store_weight_45 );
ut46_nn_multiplication: nn_multiplication port map(weight_46 , x_46 ,store_weight_46 );
ut47_nn_multiplication: nn_multiplication port map(weight_47 , x_47 ,store_weight_47 );
ut48_nn_multiplication: nn_multiplication port map(weight_48 , x_48 ,store_weight_48 );
ut49_nn_multiplication: nn_multiplication port map(weight_49 , x_49 ,store_weight_49 );
ut50_nn_multiplication: nn_multiplication port map(weight_50 , x_50 ,store_weight_50 );
ut51_nn_multiplication: nn_multiplication port map(weight_51 , x_51 ,store_weight_51 );
ut52_nn_multiplication: nn_multiplication port map(weight_52 , x_52 ,store_weight_52 );
ut53_nn_multiplication: nn_multiplication port map(weight_53 , x_53 ,store_weight_53 );
ut54_nn_multiplication: nn_multiplication port map(weight_54 , x_54 ,store_weight_54 );
ut55_nn_multiplication: nn_multiplication port map(weight_55 , x_55 ,store_weight_55 );
ut56_nn_multiplication: nn_multiplication port map(weight_56 , x_56 ,store_weight_56 );
ut57_nn_multiplication: nn_multiplication port map(weight_57 , x_57 ,store_weight_57 );
ut58_nn_multiplication: nn_multiplication port map(weight_58 , x_58 ,store_weight_58 );
ut59_nn_multiplication: nn_multiplication port map(weight_59 , x_59 ,store_weight_59 );
ut60_nn_multiplication: nn_multiplication port map(weight_60 , x_60 ,store_weight_60 );
ut61_nn_multiplication: nn_multiplication port map(weight_61 , x_61 ,store_weight_61 );
ut62_nn_multiplication: nn_multiplication port map(weight_62 , x_62 ,store_weight_62 );
ut63_nn_multiplication: nn_multiplication port map(weight_63 , x_63 ,store_weight_63 );
ut64_nn_multiplication: nn_multiplication port map(weight_64 , x_64 ,store_weight_64 );
ut65_nn_multiplication: nn_multiplication port map(weight_65 , x_65 ,store_weight_65 );
ut66_nn_multiplication: nn_multiplication port map(weight_66 , x_66 ,store_weight_66 );
ut67_nn_multiplication: nn_multiplication port map(weight_67 , x_67 ,store_weight_67 );
ut68_nn_multiplication: nn_multiplication port map(weight_68 , x_68 ,store_weight_68 );
ut69_nn_multiplication: nn_multiplication port map(weight_69 , x_69 ,store_weight_69 );
ut70_nn_multiplication: nn_multiplication port map(weight_70 , x_70 ,store_weight_70 );
ut71_nn_multiplication: nn_multiplication port map(weight_71 , x_71 ,store_weight_71 );
ut72_nn_multiplication: nn_multiplication port map(weight_72 , x_72 ,store_weight_72 );
ut73_nn_multiplication: nn_multiplication port map(weight_73 , x_73 ,store_weight_73 );
ut74_nn_multiplication: nn_multiplication port map(weight_74 , x_74 ,store_weight_74 );
ut75_nn_multiplication: nn_multiplication port map(weight_75 , x_75 ,store_weight_75 );
ut76_nn_multiplication: nn_multiplication port map(weight_76 , x_76 ,store_weight_76 );
ut77_nn_multiplication: nn_multiplication port map(weight_77 , x_77 ,store_weight_77 );
ut78_nn_multiplication: nn_multiplication port map(weight_78 , x_78 ,store_weight_78 );
ut79_nn_multiplication: nn_multiplication port map(weight_79 , x_79 ,store_weight_79 );
ut80_nn_multiplication: nn_multiplication port map(weight_80 , x_80 ,store_weight_80 );
ut81_nn_multiplication: nn_multiplication port map(weight_81 , x_81 ,store_weight_81 );
ut82_nn_multiplication: nn_multiplication port map(weight_82 , x_82 ,store_weight_82 );
ut83_nn_multiplication: nn_multiplication port map(weight_83 , x_83 ,store_weight_83 );
ut84_nn_multiplication: nn_multiplication port map(weight_84 , x_84 ,store_weight_84 );
ut85_nn_multiplication: nn_multiplication port map(weight_85 , x_85 ,store_weight_85 );
ut86_nn_multiplication: nn_multiplication port map(weight_86 , x_86 ,store_weight_86 );
ut87_nn_multiplication: nn_multiplication port map(weight_87 , x_87 ,store_weight_87 );
ut88_nn_multiplication: nn_multiplication port map(weight_88 , x_88 ,store_weight_88 );
ut89_nn_multiplication: nn_multiplication port map(weight_89 , x_89 ,store_weight_89 );
ut90_nn_multiplication: nn_multiplication port map(weight_90 , x_90 ,store_weight_90 );
ut91_nn_multiplication: nn_multiplication port map(weight_91 , x_91 ,store_weight_91 );
ut92_nn_multiplication: nn_multiplication port map(weight_92 , x_92 ,store_weight_92 );
ut93_nn_multiplication: nn_multiplication port map(weight_93 , x_93 ,store_weight_93 );
ut94_nn_multiplication: nn_multiplication port map(weight_94 , x_94 ,store_weight_94 );
ut95_nn_multiplication: nn_multiplication port map(weight_95 , x_95 ,store_weight_95 );
ut96_nn_multiplication: nn_multiplication port map(weight_96 , x_96 ,store_weight_96 );
ut97_nn_multiplication: nn_multiplication port map(weight_97 , x_97 ,store_weight_97 );
ut98_nn_multiplication: nn_multiplication port map(weight_98 , x_98 ,store_weight_98 );
ut99_nn_multiplication: nn_multiplication port map(weight_99 , x_99 ,store_weight_99 );
ut100_nn_multiplication: nn_multiplication port map(weight_100 , x_100 ,store_weight_100 );
ut101_nn_multiplication: nn_multiplication port map(weight_101 , x_101 ,store_weight_101 );
ut102_nn_multiplication: nn_multiplication port map(weight_102 , x_102 ,store_weight_102 );
ut103_nn_multiplication: nn_multiplication port map(weight_103 , x_103 ,store_weight_103 );
ut104_nn_multiplication: nn_multiplication port map(weight_104 , x_104 ,store_weight_104 );
ut105_nn_multiplication: nn_multiplication port map(weight_105 , x_105 ,store_weight_105 );
ut106_nn_multiplication: nn_multiplication port map(weight_106 , x_106 ,store_weight_106 );
ut107_nn_multiplication: nn_multiplication port map(weight_107 , x_107 ,store_weight_107 );
ut108_nn_multiplication: nn_multiplication port map(weight_108 , x_108 ,store_weight_108 );
ut109_nn_multiplication: nn_multiplication port map(weight_109 , x_109 ,store_weight_109 );
ut110_nn_multiplication: nn_multiplication port map(weight_110 , x_110 ,store_weight_110 );
ut111_nn_multiplication: nn_multiplication port map(weight_111 , x_111 ,store_weight_111 );
ut112_nn_multiplication: nn_multiplication port map(weight_112 , x_112 ,store_weight_112 );
ut113_nn_multiplication: nn_multiplication port map(weight_113 , x_113 ,store_weight_113 );
ut114_nn_multiplication: nn_multiplication port map(weight_114 , x_114 ,store_weight_114 );
ut115_nn_multiplication: nn_multiplication port map(weight_115 , x_115 ,store_weight_115 );
ut116_nn_multiplication: nn_multiplication port map(weight_116 , x_116 ,store_weight_116 );
ut117_nn_multiplication: nn_multiplication port map(weight_117 , x_117 ,store_weight_117 );
ut118_nn_multiplication: nn_multiplication port map(weight_118 , x_118 ,store_weight_118 );
ut119_nn_multiplication: nn_multiplication port map(weight_119 , x_119 ,store_weight_119 );
ut120_nn_multiplication: nn_multiplication port map(weight_120 , x_120 ,store_weight_120 );
ut121_nn_multiplication: nn_multiplication port map(weight_121 , x_121 ,store_weight_121 );
ut122_nn_multiplication: nn_multiplication port map(weight_122 , x_122 ,store_weight_122 );
ut123_nn_multiplication: nn_multiplication port map(weight_123 , x_123 ,store_weight_123 );
ut124_nn_multiplication: nn_multiplication port map(weight_124 , x_124 ,store_weight_124 );
ut125_nn_multiplication: nn_multiplication port map(weight_125 , x_125 ,store_weight_125 );
ut126_nn_multiplication: nn_multiplication port map(weight_126 , x_126 ,store_weight_126 );
ut127_nn_multiplication: nn_multiplication port map(weight_127 , x_127 ,store_weight_127 );
ut128_nn_multiplication: nn_multiplication port map(weight_128 , x_128 ,store_weight_128 );
ut129_nn_multiplication: nn_multiplication port map(weight_129 , x_129 ,store_weight_129 );
ut130_nn_multiplication: nn_multiplication port map(weight_130 , x_130 ,store_weight_130 );
ut131_nn_multiplication: nn_multiplication port map(weight_131 , x_131 ,store_weight_131 );
ut132_nn_multiplication: nn_multiplication port map(weight_132 , x_132 ,store_weight_132 );
ut133_nn_multiplication: nn_multiplication port map(weight_133 , x_133 ,store_weight_133 );
ut134_nn_multiplication: nn_multiplication port map(weight_134 , x_134 ,store_weight_134 );
ut135_nn_multiplication: nn_multiplication port map(weight_135 , x_135 ,store_weight_135 );
ut136_nn_multiplication: nn_multiplication port map(weight_136 , x_136 ,store_weight_136 );
ut137_nn_multiplication: nn_multiplication port map(weight_137 , x_137 ,store_weight_137 );
ut138_nn_multiplication: nn_multiplication port map(weight_138 , x_138 ,store_weight_138 );
ut139_nn_multiplication: nn_multiplication port map(weight_139 , x_139 ,store_weight_139 );
ut140_nn_multiplication: nn_multiplication port map(weight_140 , x_140 ,store_weight_140 );
ut141_nn_multiplication: nn_multiplication port map(weight_141 , x_141 ,store_weight_141 );
ut142_nn_multiplication: nn_multiplication port map(weight_142 , x_142 ,store_weight_142 );
ut143_nn_multiplication: nn_multiplication port map(weight_143 , x_143 ,store_weight_143 );
ut144_nn_multiplication: nn_multiplication port map(weight_144 , x_144 ,store_weight_144 );
ut145_nn_multiplication: nn_multiplication port map(weight_145 , x_145 ,store_weight_145 );
ut146_nn_multiplication: nn_multiplication port map(weight_146 , x_146 ,store_weight_146 );
ut147_nn_multiplication: nn_multiplication port map(weight_147 , x_147 ,store_weight_147 );
ut148_nn_multiplication: nn_multiplication port map(weight_148 , x_148 ,store_weight_148 );
ut149_nn_multiplication: nn_multiplication port map(weight_149 , x_149 ,store_weight_149 );
ut150_nn_multiplication: nn_multiplication port map(weight_150 , x_150 ,store_weight_150 );
ut151_nn_multiplication: nn_multiplication port map(weight_151 , x_151 ,store_weight_151 );
ut152_nn_multiplication: nn_multiplication port map(weight_152 , x_152 ,store_weight_152 );
ut153_nn_multiplication: nn_multiplication port map(weight_153 , x_153 ,store_weight_153 );
ut154_nn_multiplication: nn_multiplication port map(weight_154 , x_154 ,store_weight_154 );
ut155_nn_multiplication: nn_multiplication port map(weight_155 , x_155 ,store_weight_155 );
ut156_nn_multiplication: nn_multiplication port map(weight_156 , x_156 ,store_weight_156 );
ut157_nn_multiplication: nn_multiplication port map(weight_157 , x_157 ,store_weight_157 );
ut158_nn_multiplication: nn_multiplication port map(weight_158 , x_158 ,store_weight_158 );
ut159_nn_multiplication: nn_multiplication port map(weight_159 , x_159 ,store_weight_159 );
ut160_nn_multiplication: nn_multiplication port map(weight_160 , x_160 ,store_weight_160 );
ut161_nn_multiplication: nn_multiplication port map(weight_161 , x_161 ,store_weight_161 );
ut162_nn_multiplication: nn_multiplication port map(weight_162 , x_162 ,store_weight_162 );
ut163_nn_multiplication: nn_multiplication port map(weight_163 , x_163 ,store_weight_163 );
ut164_nn_multiplication: nn_multiplication port map(weight_164 , x_164 ,store_weight_164 );
ut165_nn_multiplication: nn_multiplication port map(weight_165 , x_165 ,store_weight_165 );
ut166_nn_multiplication: nn_multiplication port map(weight_166 , x_166 ,store_weight_166 );
ut167_nn_multiplication: nn_multiplication port map(weight_167 , x_167 ,store_weight_167 );
ut168_nn_multiplication: nn_multiplication port map(weight_168 , x_168 ,store_weight_168 );
ut169_nn_multiplication: nn_multiplication port map(weight_169 , x_169 ,store_weight_169 );
ut170_nn_multiplication: nn_multiplication port map(weight_170 , x_170 ,store_weight_170 );
ut171_nn_multiplication: nn_multiplication port map(weight_171 , x_171 ,store_weight_171 );
ut172_nn_multiplication: nn_multiplication port map(weight_172 , x_172 ,store_weight_172 );
ut173_nn_multiplication: nn_multiplication port map(weight_173 , x_173 ,store_weight_173 );
ut174_nn_multiplication: nn_multiplication port map(weight_174 , x_174 ,store_weight_174 );
ut175_nn_multiplication: nn_multiplication port map(weight_175 , x_175 ,store_weight_175 );
ut176_nn_multiplication: nn_multiplication port map(weight_176 , x_176 ,store_weight_176 );
ut177_nn_multiplication: nn_multiplication port map(weight_177 , x_177 ,store_weight_177 );
ut178_nn_multiplication: nn_multiplication port map(weight_178 , x_178 ,store_weight_178 );
ut179_nn_multiplication: nn_multiplication port map(weight_179 , x_179 ,store_weight_179 );
ut180_nn_multiplication: nn_multiplication port map(weight_180 , x_180 ,store_weight_180 );
ut181_nn_multiplication: nn_multiplication port map(weight_181 , x_181 ,store_weight_181 );
ut182_nn_multiplication: nn_multiplication port map(weight_182 , x_182 ,store_weight_182 );
ut183_nn_multiplication: nn_multiplication port map(weight_183 , x_183 ,store_weight_183 );
ut184_nn_multiplication: nn_multiplication port map(weight_184 , x_184 ,store_weight_184 );
ut185_nn_multiplication: nn_multiplication port map(weight_185 , x_185 ,store_weight_185 );
ut186_nn_multiplication: nn_multiplication port map(weight_186 , x_186 ,store_weight_186 );
ut187_nn_multiplication: nn_multiplication port map(weight_187 , x_187 ,store_weight_187 );
ut188_nn_multiplication: nn_multiplication port map(weight_188 , x_188 ,store_weight_188 );
ut189_nn_multiplication: nn_multiplication port map(weight_189 , x_189 ,store_weight_189 );
ut190_nn_multiplication: nn_multiplication port map(weight_190 , x_190 ,store_weight_190 );
ut191_nn_multiplication: nn_multiplication port map(weight_191 , x_191 ,store_weight_191 );
ut192_nn_multiplication: nn_multiplication port map(weight_192 , x_192 ,store_weight_192 );
ut193_nn_multiplication: nn_multiplication port map(weight_193 , x_193 ,store_weight_193 );
ut194_nn_multiplication: nn_multiplication port map(weight_194 , x_194 ,store_weight_194 );
ut195_nn_multiplication: nn_multiplication port map(weight_195 , x_195 ,store_weight_195 );
ut196_nn_multiplication: nn_multiplication port map(weight_196 , x_196 ,store_weight_196 );
ut197_nn_multiplication: nn_multiplication port map(weight_197 , x_197 ,store_weight_197 );
ut198_nn_multiplication: nn_multiplication port map(weight_198 , x_198 ,store_weight_198 );
ut199_nn_multiplication: nn_multiplication port map(weight_199 , x_199 ,store_weight_199 );
ut200_nn_multiplication: nn_multiplication port map(weight_200 , x_200 ,store_weight_200 );
ut201_nn_multiplication: nn_multiplication port map(weight_201 , x_201 ,store_weight_201 );
ut202_nn_multiplication: nn_multiplication port map(weight_202 , x_202 ,store_weight_202 );
ut203_nn_multiplication: nn_multiplication port map(weight_203 , x_203 ,store_weight_203 );
ut204_nn_multiplication: nn_multiplication port map(weight_204 , x_204 ,store_weight_204 );
ut205_nn_multiplication: nn_multiplication port map(weight_205 , x_205 ,store_weight_205 );
ut206_nn_multiplication: nn_multiplication port map(weight_206 , x_206 ,store_weight_206 );
ut207_nn_multiplication: nn_multiplication port map(weight_207 , x_207 ,store_weight_207 );
ut208_nn_multiplication: nn_multiplication port map(weight_208 , x_208 ,store_weight_208 );
ut209_nn_multiplication: nn_multiplication port map(weight_209 , x_209 ,store_weight_209 );
ut210_nn_multiplication: nn_multiplication port map(weight_210 , x_210 ,store_weight_210 );
ut211_nn_multiplication: nn_multiplication port map(weight_211 , x_211 ,store_weight_211 );
ut212_nn_multiplication: nn_multiplication port map(weight_212 , x_212 ,store_weight_212 );
ut213_nn_multiplication: nn_multiplication port map(weight_213 , x_213 ,store_weight_213 );
ut214_nn_multiplication: nn_multiplication port map(weight_214 , x_214 ,store_weight_214 );
ut215_nn_multiplication: nn_multiplication port map(weight_215 , x_215 ,store_weight_215 );
ut216_nn_multiplication: nn_multiplication port map(weight_216 , x_216 ,store_weight_216 );
ut217_nn_multiplication: nn_multiplication port map(weight_217 , x_217 ,store_weight_217 );
ut218_nn_multiplication: nn_multiplication port map(weight_218 , x_218 ,store_weight_218 );
ut219_nn_multiplication: nn_multiplication port map(weight_219 , x_219 ,store_weight_219 );
ut220_nn_multiplication: nn_multiplication port map(weight_220 , x_220 ,store_weight_220 );
ut221_nn_multiplication: nn_multiplication port map(weight_221 , x_221 ,store_weight_221 );
ut222_nn_multiplication: nn_multiplication port map(weight_222 , x_222 ,store_weight_222 );
ut223_nn_multiplication: nn_multiplication port map(weight_223 , x_223 ,store_weight_223 );
ut224_nn_multiplication: nn_multiplication port map(weight_224 , x_224 ,store_weight_224 );
ut225_nn_multiplication: nn_multiplication port map(weight_225 , x_225 ,store_weight_225 );
ut226_nn_multiplication: nn_multiplication port map(weight_226 , x_226 ,store_weight_226 );
ut227_nn_multiplication: nn_multiplication port map(weight_227 , x_227 ,store_weight_227 );
ut228_nn_multiplication: nn_multiplication port map(weight_228 , x_228 ,store_weight_228 );
ut229_nn_multiplication: nn_multiplication port map(weight_229 , x_229 ,store_weight_229 );
ut230_nn_multiplication: nn_multiplication port map(weight_230 , x_230 ,store_weight_230 );
ut231_nn_multiplication: nn_multiplication port map(weight_231 , x_231 ,store_weight_231 );
ut232_nn_multiplication: nn_multiplication port map(weight_232 , x_232 ,store_weight_232 );
ut233_nn_multiplication: nn_multiplication port map(weight_233 , x_233 ,store_weight_233 );
ut234_nn_multiplication: nn_multiplication port map(weight_234 , x_234 ,store_weight_234 );
ut235_nn_multiplication: nn_multiplication port map(weight_235 , x_235 ,store_weight_235 );
ut236_nn_multiplication: nn_multiplication port map(weight_236 , x_236 ,store_weight_236 );
ut237_nn_multiplication: nn_multiplication port map(weight_237 , x_237 ,store_weight_237 );
ut238_nn_multiplication: nn_multiplication port map(weight_238 , x_238 ,store_weight_238 );
ut239_nn_multiplication: nn_multiplication port map(weight_239 , x_239 ,store_weight_239 );
ut240_nn_multiplication: nn_multiplication port map(weight_240 , x_240 ,store_weight_240 );
ut241_nn_multiplication: nn_multiplication port map(weight_241 , x_241 ,store_weight_241 );
ut242_nn_multiplication: nn_multiplication port map(weight_242 , x_242 ,store_weight_242 );
ut243_nn_multiplication: nn_multiplication port map(weight_243 , x_243 ,store_weight_243 );
ut244_nn_multiplication: nn_multiplication port map(weight_244 , x_244 ,store_weight_244 );
ut245_nn_multiplication: nn_multiplication port map(weight_245 , x_245 ,store_weight_245 );
ut246_nn_multiplication: nn_multiplication port map(weight_246 , x_246 ,store_weight_246 );
ut247_nn_multiplication: nn_multiplication port map(weight_247 , x_247 ,store_weight_247 );
ut248_nn_multiplication: nn_multiplication port map(weight_248 , x_248 ,store_weight_248 );
ut249_nn_multiplication: nn_multiplication port map(weight_249 , x_249 ,store_weight_249 );
ut250_nn_multiplication: nn_multiplication port map(weight_250 , x_250 ,store_weight_250 );
ut251_nn_multiplication: nn_multiplication port map(weight_251 , x_251 ,store_weight_251 );
ut252_nn_multiplication: nn_multiplication port map(weight_252 , x_252 ,store_weight_252 );
ut253_nn_multiplication: nn_multiplication port map(weight_253 , x_253 ,store_weight_253 );
ut254_nn_multiplication: nn_multiplication port map(weight_254 , x_254 ,store_weight_254 );
ut255_nn_multiplication: nn_multiplication port map(weight_255 , x_255 ,store_weight_255 );
ut256_nn_multiplication: nn_multiplication port map(weight_256 , x_256 ,store_weight_256 );
ut257_nn_multiplication: nn_multiplication port map(weight_257 , x_257 ,store_weight_257 );
ut258_nn_multiplication: nn_multiplication port map(weight_258 , x_258 ,store_weight_258 );
ut259_nn_multiplication: nn_multiplication port map(weight_259 , x_259 ,store_weight_259 );
ut260_nn_multiplication: nn_multiplication port map(weight_260 , x_260 ,store_weight_260 );
ut261_nn_multiplication: nn_multiplication port map(weight_261 , x_261 ,store_weight_261 );
ut262_nn_multiplication: nn_multiplication port map(weight_262 , x_262 ,store_weight_262 );
ut263_nn_multiplication: nn_multiplication port map(weight_263 , x_263 ,store_weight_263 );
ut264_nn_multiplication: nn_multiplication port map(weight_264 , x_264 ,store_weight_264 );
ut265_nn_multiplication: nn_multiplication port map(weight_265 , x_265 ,store_weight_265 );
ut266_nn_multiplication: nn_multiplication port map(weight_266 , x_266 ,store_weight_266 );
ut267_nn_multiplication: nn_multiplication port map(weight_267 , x_267 ,store_weight_267 );
ut268_nn_multiplication: nn_multiplication port map(weight_268 , x_268 ,store_weight_268 );
ut269_nn_multiplication: nn_multiplication port map(weight_269 , x_269 ,store_weight_269 );
ut270_nn_multiplication: nn_multiplication port map(weight_270 , x_270 ,store_weight_270 );
ut271_nn_multiplication: nn_multiplication port map(weight_271 , x_271 ,store_weight_271 );
ut272_nn_multiplication: nn_multiplication port map(weight_272 , x_272 ,store_weight_272 );
ut273_nn_multiplication: nn_multiplication port map(weight_273 , x_273 ,store_weight_273 );
ut274_nn_multiplication: nn_multiplication port map(weight_274 , x_274 ,store_weight_274 );
ut275_nn_multiplication: nn_multiplication port map(weight_275 , x_275 ,store_weight_275 );
ut276_nn_multiplication: nn_multiplication port map(weight_276 , x_276 ,store_weight_276 );
ut277_nn_multiplication: nn_multiplication port map(weight_277 , x_277 ,store_weight_277 );
ut278_nn_multiplication: nn_multiplication port map(weight_278 , x_278 ,store_weight_278 );
ut279_nn_multiplication: nn_multiplication port map(weight_279 , x_279 ,store_weight_279 );
ut280_nn_multiplication: nn_multiplication port map(weight_280 , x_280 ,store_weight_280 );
ut281_nn_multiplication: nn_multiplication port map(weight_281 , x_281 ,store_weight_281 );
ut282_nn_multiplication: nn_multiplication port map(weight_282 , x_282 ,store_weight_282 );
ut283_nn_multiplication: nn_multiplication port map(weight_283 , x_283 ,store_weight_283 );
ut284_nn_multiplication: nn_multiplication port map(weight_284 , x_284 ,store_weight_284 );
ut285_nn_multiplication: nn_multiplication port map(weight_285 , x_285 ,store_weight_285 );
ut286_nn_multiplication: nn_multiplication port map(weight_286 , x_286 ,store_weight_286 );
ut287_nn_multiplication: nn_multiplication port map(weight_287 , x_287 ,store_weight_287 );
ut288_nn_multiplication: nn_multiplication port map(weight_288 , x_288 ,store_weight_288 );
ut289_nn_multiplication: nn_multiplication port map(weight_289 , x_289 ,store_weight_289 );
ut290_nn_multiplication: nn_multiplication port map(weight_290 , x_290 ,store_weight_290 );
ut291_nn_multiplication: nn_multiplication port map(weight_291 , x_291 ,store_weight_291 );
ut292_nn_multiplication: nn_multiplication port map(weight_292 , x_292 ,store_weight_292 );
ut293_nn_multiplication: nn_multiplication port map(weight_293 , x_293 ,store_weight_293 );
ut294_nn_multiplication: nn_multiplication port map(weight_294 , x_294 ,store_weight_294 );
ut295_nn_multiplication: nn_multiplication port map(weight_295 , x_295 ,store_weight_295 );
ut296_nn_multiplication: nn_multiplication port map(weight_296 , x_296 ,store_weight_296 );
ut297_nn_multiplication: nn_multiplication port map(weight_297 , x_297 ,store_weight_297 );
ut298_nn_multiplication: nn_multiplication port map(weight_298 , x_298 ,store_weight_298 );
ut299_nn_multiplication: nn_multiplication port map(weight_299 , x_299 ,store_weight_299 );
ut300_nn_multiplication: nn_multiplication port map(weight_300 , x_300 ,store_weight_300 );
ut301_nn_multiplication: nn_multiplication port map(weight_301 , x_301 ,store_weight_301 );
ut302_nn_multiplication: nn_multiplication port map(weight_302 , x_302 ,store_weight_302 );
ut303_nn_multiplication: nn_multiplication port map(weight_303 , x_303 ,store_weight_303 );
ut304_nn_multiplication: nn_multiplication port map(weight_304 , x_304 ,store_weight_304 );
ut305_nn_multiplication: nn_multiplication port map(weight_305 , x_305 ,store_weight_305 );
ut306_nn_multiplication: nn_multiplication port map(weight_306 , x_306 ,store_weight_306 );
ut307_nn_multiplication: nn_multiplication port map(weight_307 , x_307 ,store_weight_307 );
ut308_nn_multiplication: nn_multiplication port map(weight_308 , x_308 ,store_weight_308 );
ut309_nn_multiplication: nn_multiplication port map(weight_309 , x_309 ,store_weight_309 );
ut310_nn_multiplication: nn_multiplication port map(weight_310 , x_310 ,store_weight_310 );
ut311_nn_multiplication: nn_multiplication port map(weight_311 , x_311 ,store_weight_311 );
ut312_nn_multiplication: nn_multiplication port map(weight_312 , x_312 ,store_weight_312 );
ut313_nn_multiplication: nn_multiplication port map(weight_313 , x_313 ,store_weight_313 );
ut314_nn_multiplication: nn_multiplication port map(weight_314 , x_314 ,store_weight_314 );
ut315_nn_multiplication: nn_multiplication port map(weight_315 , x_315 ,store_weight_315 );
ut316_nn_multiplication: nn_multiplication port map(weight_316 , x_316 ,store_weight_316 );
ut317_nn_multiplication: nn_multiplication port map(weight_317 , x_317 ,store_weight_317 );
ut318_nn_multiplication: nn_multiplication port map(weight_318 , x_318 ,store_weight_318 );
ut319_nn_multiplication: nn_multiplication port map(weight_319 , x_319 ,store_weight_319 );
ut320_nn_multiplication: nn_multiplication port map(weight_320 , x_320 ,store_weight_320 );
ut321_nn_multiplication: nn_multiplication port map(weight_321 , x_321 ,store_weight_321 );
ut322_nn_multiplication: nn_multiplication port map(weight_322 , x_322 ,store_weight_322 );
ut323_nn_multiplication: nn_multiplication port map(weight_323 , x_323 ,store_weight_323 );
ut324_nn_multiplication: nn_multiplication port map(weight_324 , x_324 ,store_weight_324 );
ut325_nn_multiplication: nn_multiplication port map(weight_325 , x_325 ,store_weight_325 );
ut326_nn_multiplication: nn_multiplication port map(weight_326 , x_326 ,store_weight_326 );
ut327_nn_multiplication: nn_multiplication port map(weight_327 , x_327 ,store_weight_327 );
ut328_nn_multiplication: nn_multiplication port map(weight_328 , x_328 ,store_weight_328 );
ut329_nn_multiplication: nn_multiplication port map(weight_329 , x_329 ,store_weight_329 );
ut330_nn_multiplication: nn_multiplication port map(weight_330 , x_330 ,store_weight_330 );
ut331_nn_multiplication: nn_multiplication port map(weight_331 , x_331 ,store_weight_331 );
ut332_nn_multiplication: nn_multiplication port map(weight_332 , x_332 ,store_weight_332 );
ut333_nn_multiplication: nn_multiplication port map(weight_333 , x_333 ,store_weight_333 );
ut334_nn_multiplication: nn_multiplication port map(weight_334 , x_334 ,store_weight_334 );
ut335_nn_multiplication: nn_multiplication port map(weight_335 , x_335 ,store_weight_335 );
ut336_nn_multiplication: nn_multiplication port map(weight_336 , x_336 ,store_weight_336 );
ut337_nn_multiplication: nn_multiplication port map(weight_337 , x_337 ,store_weight_337 );
ut338_nn_multiplication: nn_multiplication port map(weight_338 , x_338 ,store_weight_338 );
ut339_nn_multiplication: nn_multiplication port map(weight_339 , x_339 ,store_weight_339 );
ut340_nn_multiplication: nn_multiplication port map(weight_340 , x_340 ,store_weight_340 );
ut341_nn_multiplication: nn_multiplication port map(weight_341 , x_341 ,store_weight_341 );
ut342_nn_multiplication: nn_multiplication port map(weight_342 , x_342 ,store_weight_342 );
ut343_nn_multiplication: nn_multiplication port map(weight_343 , x_343 ,store_weight_343 );
ut344_nn_multiplication: nn_multiplication port map(weight_344 , x_344 ,store_weight_344 );
ut345_nn_multiplication: nn_multiplication port map(weight_345 , x_345 ,store_weight_345 );
ut346_nn_multiplication: nn_multiplication port map(weight_346 , x_346 ,store_weight_346 );
ut347_nn_multiplication: nn_multiplication port map(weight_347 , x_347 ,store_weight_347 );
ut348_nn_multiplication: nn_multiplication port map(weight_348 , x_348 ,store_weight_348 );
ut349_nn_multiplication: nn_multiplication port map(weight_349 , x_349 ,store_weight_349 );
ut350_nn_multiplication: nn_multiplication port map(weight_350 , x_350 ,store_weight_350 );
ut351_nn_multiplication: nn_multiplication port map(weight_351 , x_351 ,store_weight_351 );
ut352_nn_multiplication: nn_multiplication port map(weight_352 , x_352 ,store_weight_352 );
ut353_nn_multiplication: nn_multiplication port map(weight_353 , x_353 ,store_weight_353 );
ut354_nn_multiplication: nn_multiplication port map(weight_354 , x_354 ,store_weight_354 );
ut355_nn_multiplication: nn_multiplication port map(weight_355 , x_355 ,store_weight_355 );
ut356_nn_multiplication: nn_multiplication port map(weight_356 , x_356 ,store_weight_356 );
ut357_nn_multiplication: nn_multiplication port map(weight_357 , x_357 ,store_weight_357 );
ut358_nn_multiplication: nn_multiplication port map(weight_358 , x_358 ,store_weight_358 );
ut359_nn_multiplication: nn_multiplication port map(weight_359 , x_359 ,store_weight_359 );
ut360_nn_multiplication: nn_multiplication port map(weight_360 , x_360 ,store_weight_360 );
ut361_nn_multiplication: nn_multiplication port map(weight_361 , x_361 ,store_weight_361 );
ut362_nn_multiplication: nn_multiplication port map(weight_362 , x_362 ,store_weight_362 );
ut363_nn_multiplication: nn_multiplication port map(weight_363 , x_363 ,store_weight_363 );
ut364_nn_multiplication: nn_multiplication port map(weight_364 , x_364 ,store_weight_364 );
ut365_nn_multiplication: nn_multiplication port map(weight_365 , x_365 ,store_weight_365 );
ut366_nn_multiplication: nn_multiplication port map(weight_366 , x_366 ,store_weight_366 );
ut367_nn_multiplication: nn_multiplication port map(weight_367 , x_367 ,store_weight_367 );
ut368_nn_multiplication: nn_multiplication port map(weight_368 , x_368 ,store_weight_368 );
ut369_nn_multiplication: nn_multiplication port map(weight_369 , x_369 ,store_weight_369 );
ut370_nn_multiplication: nn_multiplication port map(weight_370 , x_370 ,store_weight_370 );
ut371_nn_multiplication: nn_multiplication port map(weight_371 , x_371 ,store_weight_371 );
ut372_nn_multiplication: nn_multiplication port map(weight_372 , x_372 ,store_weight_372 );
ut373_nn_multiplication: nn_multiplication port map(weight_373 , x_373 ,store_weight_373 );
ut374_nn_multiplication: nn_multiplication port map(weight_374 , x_374 ,store_weight_374 );
ut375_nn_multiplication: nn_multiplication port map(weight_375 , x_375 ,store_weight_375 );
ut376_nn_multiplication: nn_multiplication port map(weight_376 , x_376 ,store_weight_376 );
ut377_nn_multiplication: nn_multiplication port map(weight_377 , x_377 ,store_weight_377 );
ut378_nn_multiplication: nn_multiplication port map(weight_378 , x_378 ,store_weight_378 );
ut379_nn_multiplication: nn_multiplication port map(weight_379 , x_379 ,store_weight_379 );
ut380_nn_multiplication: nn_multiplication port map(weight_380 , x_380 ,store_weight_380 );
ut381_nn_multiplication: nn_multiplication port map(weight_381 , x_381 ,store_weight_381 );
ut382_nn_multiplication: nn_multiplication port map(weight_382 , x_382 ,store_weight_382 );
ut383_nn_multiplication: nn_multiplication port map(weight_383 , x_383 ,store_weight_383 );
ut384_nn_multiplication: nn_multiplication port map(weight_384 , x_384 ,store_weight_384 );
ut385_nn_multiplication: nn_multiplication port map(weight_385 , x_385 ,store_weight_385 );
ut386_nn_multiplication: nn_multiplication port map(weight_386 , x_386 ,store_weight_386 );
ut387_nn_multiplication: nn_multiplication port map(weight_387 , x_387 ,store_weight_387 );
ut388_nn_multiplication: nn_multiplication port map(weight_388 , x_388 ,store_weight_388 );
ut389_nn_multiplication: nn_multiplication port map(weight_389 , x_389 ,store_weight_389 );
ut390_nn_multiplication: nn_multiplication port map(weight_390 , x_390 ,store_weight_390 );
ut391_nn_multiplication: nn_multiplication port map(weight_391 , x_391 ,store_weight_391 );
ut392_nn_multiplication: nn_multiplication port map(weight_392 , x_392 ,store_weight_392 );
ut393_nn_multiplication: nn_multiplication port map(weight_393 , x_393 ,store_weight_393 );
ut394_nn_multiplication: nn_multiplication port map(weight_394 , x_394 ,store_weight_394 );
ut395_nn_multiplication: nn_multiplication port map(weight_395 , x_395 ,store_weight_395 );
ut396_nn_multiplication: nn_multiplication port map(weight_396 , x_396 ,store_weight_396 );
ut397_nn_multiplication: nn_multiplication port map(weight_397 , x_397 ,store_weight_397 );
ut398_nn_multiplication: nn_multiplication port map(weight_398 , x_398 ,store_weight_398 );
ut399_nn_multiplication: nn_multiplication port map(weight_399 , x_399 ,store_weight_399 );
ut400_nn_multiplication: nn_multiplication port map(weight_400 , x_400 ,store_weight_400 );
ut401_nn_multiplication: nn_multiplication port map(weight_401 , x_401 ,store_weight_401 );
ut402_nn_multiplication: nn_multiplication port map(weight_402 , x_402 ,store_weight_402 );
ut403_nn_multiplication: nn_multiplication port map(weight_403 , x_403 ,store_weight_403 );
ut404_nn_multiplication: nn_multiplication port map(weight_404 , x_404 ,store_weight_404 );
ut405_nn_multiplication: nn_multiplication port map(weight_405 , x_405 ,store_weight_405 );
ut406_nn_multiplication: nn_multiplication port map(weight_406 , x_406 ,store_weight_406 );
ut407_nn_multiplication: nn_multiplication port map(weight_407 , x_407 ,store_weight_407 );
ut408_nn_multiplication: nn_multiplication port map(weight_408 , x_408 ,store_weight_408 );
ut409_nn_multiplication: nn_multiplication port map(weight_409 , x_409 ,store_weight_409 );
ut410_nn_multiplication: nn_multiplication port map(weight_410 , x_410 ,store_weight_410 );
ut411_nn_multiplication: nn_multiplication port map(weight_411 , x_411 ,store_weight_411 );
ut412_nn_multiplication: nn_multiplication port map(weight_412 , x_412 ,store_weight_412 );
ut413_nn_multiplication: nn_multiplication port map(weight_413 , x_413 ,store_weight_413 );
ut414_nn_multiplication: nn_multiplication port map(weight_414 , x_414 ,store_weight_414 );
ut415_nn_multiplication: nn_multiplication port map(weight_415 , x_415 ,store_weight_415 );
ut416_nn_multiplication: nn_multiplication port map(weight_416 , x_416 ,store_weight_416 );
ut417_nn_multiplication: nn_multiplication port map(weight_417 , x_417 ,store_weight_417 );
ut418_nn_multiplication: nn_multiplication port map(weight_418 , x_418 ,store_weight_418 );
ut419_nn_multiplication: nn_multiplication port map(weight_419 , x_419 ,store_weight_419 );
ut420_nn_multiplication: nn_multiplication port map(weight_420 , x_420 ,store_weight_420 );
ut421_nn_multiplication: nn_multiplication port map(weight_421 , x_421 ,store_weight_421 );
ut422_nn_multiplication: nn_multiplication port map(weight_422 , x_422 ,store_weight_422 );
ut423_nn_multiplication: nn_multiplication port map(weight_423 , x_423 ,store_weight_423 );
ut424_nn_multiplication: nn_multiplication port map(weight_424 , x_424 ,store_weight_424 );
ut425_nn_multiplication: nn_multiplication port map(weight_425 , x_425 ,store_weight_425 );
ut426_nn_multiplication: nn_multiplication port map(weight_426 , x_426 ,store_weight_426 );
ut427_nn_multiplication: nn_multiplication port map(weight_427 , x_427 ,store_weight_427 );
ut428_nn_multiplication: nn_multiplication port map(weight_428 , x_428 ,store_weight_428 );
ut429_nn_multiplication: nn_multiplication port map(weight_429 , x_429 ,store_weight_429 );
ut430_nn_multiplication: nn_multiplication port map(weight_430 , x_430 ,store_weight_430 );
ut431_nn_multiplication: nn_multiplication port map(weight_431 , x_431 ,store_weight_431 );
ut432_nn_multiplication: nn_multiplication port map(weight_432 , x_432 ,store_weight_432 );
ut433_nn_multiplication: nn_multiplication port map(weight_433 , x_433 ,store_weight_433 );
ut434_nn_multiplication: nn_multiplication port map(weight_434 , x_434 ,store_weight_434 );
ut435_nn_multiplication: nn_multiplication port map(weight_435 , x_435 ,store_weight_435 );
ut436_nn_multiplication: nn_multiplication port map(weight_436 , x_436 ,store_weight_436 );
ut437_nn_multiplication: nn_multiplication port map(weight_437 , x_437 ,store_weight_437 );
ut438_nn_multiplication: nn_multiplication port map(weight_438 , x_438 ,store_weight_438 );
ut439_nn_multiplication: nn_multiplication port map(weight_439 , x_439 ,store_weight_439 );
ut440_nn_multiplication: nn_multiplication port map(weight_440 , x_440 ,store_weight_440 );
ut441_nn_multiplication: nn_multiplication port map(weight_441 , x_441 ,store_weight_441 );
ut442_nn_multiplication: nn_multiplication port map(weight_442 , x_442 ,store_weight_442 );
ut443_nn_multiplication: nn_multiplication port map(weight_443 , x_443 ,store_weight_443 );
ut444_nn_multiplication: nn_multiplication port map(weight_444 , x_444 ,store_weight_444 );
ut445_nn_multiplication: nn_multiplication port map(weight_445 , x_445 ,store_weight_445 );
ut446_nn_multiplication: nn_multiplication port map(weight_446 , x_446 ,store_weight_446 );
ut447_nn_multiplication: nn_multiplication port map(weight_447 , x_447 ,store_weight_447 );
ut448_nn_multiplication: nn_multiplication port map(weight_448 , x_448 ,store_weight_448 );
ut449_nn_multiplication: nn_multiplication port map(weight_449 , x_449 ,store_weight_449 );
ut450_nn_multiplication: nn_multiplication port map(weight_450 , x_450 ,store_weight_450 );
ut451_nn_multiplication: nn_multiplication port map(weight_451 , x_451 ,store_weight_451 );
ut452_nn_multiplication: nn_multiplication port map(weight_452 , x_452 ,store_weight_452 );
ut453_nn_multiplication: nn_multiplication port map(weight_453 , x_453 ,store_weight_453 );
ut454_nn_multiplication: nn_multiplication port map(weight_454 , x_454 ,store_weight_454 );
ut455_nn_multiplication: nn_multiplication port map(weight_455 , x_455 ,store_weight_455 );
ut456_nn_multiplication: nn_multiplication port map(weight_456 , x_456 ,store_weight_456 );
ut457_nn_multiplication: nn_multiplication port map(weight_457 , x_457 ,store_weight_457 );
ut458_nn_multiplication: nn_multiplication port map(weight_458 , x_458 ,store_weight_458 );
ut459_nn_multiplication: nn_multiplication port map(weight_459 , x_459 ,store_weight_459 );
ut460_nn_multiplication: nn_multiplication port map(weight_460 , x_460 ,store_weight_460 );
ut461_nn_multiplication: nn_multiplication port map(weight_461 , x_461 ,store_weight_461 );
ut462_nn_multiplication: nn_multiplication port map(weight_462 , x_462 ,store_weight_462 );
ut463_nn_multiplication: nn_multiplication port map(weight_463 , x_463 ,store_weight_463 );
ut464_nn_multiplication: nn_multiplication port map(weight_464 , x_464 ,store_weight_464 );
ut465_nn_multiplication: nn_multiplication port map(weight_465 , x_465 ,store_weight_465 );
ut466_nn_multiplication: nn_multiplication port map(weight_466 , x_466 ,store_weight_466 );
ut467_nn_multiplication: nn_multiplication port map(weight_467 , x_467 ,store_weight_467 );
ut468_nn_multiplication: nn_multiplication port map(weight_468 , x_468 ,store_weight_468 );
ut469_nn_multiplication: nn_multiplication port map(weight_469 , x_469 ,store_weight_469 );
ut470_nn_multiplication: nn_multiplication port map(weight_470 , x_470 ,store_weight_470 );
ut471_nn_multiplication: nn_multiplication port map(weight_471 , x_471 ,store_weight_471 );
ut472_nn_multiplication: nn_multiplication port map(weight_472 , x_472 ,store_weight_472 );
ut473_nn_multiplication: nn_multiplication port map(weight_473 , x_473 ,store_weight_473 );
ut474_nn_multiplication: nn_multiplication port map(weight_474 , x_474 ,store_weight_474 );
ut475_nn_multiplication: nn_multiplication port map(weight_475 , x_475 ,store_weight_475 );
ut476_nn_multiplication: nn_multiplication port map(weight_476 , x_476 ,store_weight_476 );
ut477_nn_multiplication: nn_multiplication port map(weight_477 , x_477 ,store_weight_477 );
ut478_nn_multiplication: nn_multiplication port map(weight_478 , x_478 ,store_weight_478 );
ut479_nn_multiplication: nn_multiplication port map(weight_479 , x_479 ,store_weight_479 );
ut480_nn_multiplication: nn_multiplication port map(weight_480 , x_480 ,store_weight_480 );
ut481_nn_multiplication: nn_multiplication port map(weight_481 , x_481 ,store_weight_481 );
ut482_nn_multiplication: nn_multiplication port map(weight_482 , x_482 ,store_weight_482 );
ut483_nn_multiplication: nn_multiplication port map(weight_483 , x_483 ,store_weight_483 );
ut484_nn_multiplication: nn_multiplication port map(weight_484 , x_484 ,store_weight_484 );
ut485_nn_multiplication: nn_multiplication port map(weight_485 , x_485 ,store_weight_485 );
ut486_nn_multiplication: nn_multiplication port map(weight_486 , x_486 ,store_weight_486 );
ut487_nn_multiplication: nn_multiplication port map(weight_487 , x_487 ,store_weight_487 );
ut488_nn_multiplication: nn_multiplication port map(weight_488 , x_488 ,store_weight_488 );
ut489_nn_multiplication: nn_multiplication port map(weight_489 , x_489 ,store_weight_489 );
ut490_nn_multiplication: nn_multiplication port map(weight_490 , x_490 ,store_weight_490 );
ut491_nn_multiplication: nn_multiplication port map(weight_491 , x_491 ,store_weight_491 );
ut492_nn_multiplication: nn_multiplication port map(weight_492 , x_492 ,store_weight_492 );
ut493_nn_multiplication: nn_multiplication port map(weight_493 , x_493 ,store_weight_493 );
ut494_nn_multiplication: nn_multiplication port map(weight_494 , x_494 ,store_weight_494 );
ut495_nn_multiplication: nn_multiplication port map(weight_495 , x_495 ,store_weight_495 );
ut496_nn_multiplication: nn_multiplication port map(weight_496 , x_496 ,store_weight_496 );
ut497_nn_multiplication: nn_multiplication port map(weight_497 , x_497 ,store_weight_497 );
ut498_nn_multiplication: nn_multiplication port map(weight_498 , x_498 ,store_weight_498 );
ut499_nn_multiplication: nn_multiplication port map(weight_499 , x_499 ,store_weight_499 );
ut500_nn_multiplication: nn_multiplication port map(weight_500 , x_500 ,store_weight_500 );
ut501_nn_multiplication: nn_multiplication port map(weight_501 , x_501 ,store_weight_501 );
ut502_nn_multiplication: nn_multiplication port map(weight_502 , x_502 ,store_weight_502 );
ut503_nn_multiplication: nn_multiplication port map(weight_503 , x_503 ,store_weight_503 );
ut504_nn_multiplication: nn_multiplication port map(weight_504 , x_504 ,store_weight_504 );
ut505_nn_multiplication: nn_multiplication port map(weight_505 , x_505 ,store_weight_505 );
ut506_nn_multiplication: nn_multiplication port map(weight_506 , x_506 ,store_weight_506 );
ut507_nn_multiplication: nn_multiplication port map(weight_507 , x_507 ,store_weight_507 );
ut508_nn_multiplication: nn_multiplication port map(weight_508 , x_508 ,store_weight_508 );
ut509_nn_multiplication: nn_multiplication port map(weight_509 , x_509 ,store_weight_509 );
ut510_nn_multiplication: nn_multiplication port map(weight_510 , x_510 ,store_weight_510 );
ut511_nn_multiplication: nn_multiplication port map(weight_511 , x_511 ,store_weight_511 );
ut512_nn_multiplication: nn_multiplication port map(weight_512 , x_512 ,store_weight_512 );
ut513_nn_multiplication: nn_multiplication port map(weight_513 , x_513 ,store_weight_513 );
ut514_nn_multiplication: nn_multiplication port map(weight_514 , x_514 ,store_weight_514 );
ut515_nn_multiplication: nn_multiplication port map(weight_515 , x_515 ,store_weight_515 );
ut516_nn_multiplication: nn_multiplication port map(weight_516 , x_516 ,store_weight_516 );
ut517_nn_multiplication: nn_multiplication port map(weight_517 , x_517 ,store_weight_517 );
ut518_nn_multiplication: nn_multiplication port map(weight_518 , x_518 ,store_weight_518 );
ut519_nn_multiplication: nn_multiplication port map(weight_519 , x_519 ,store_weight_519 );
ut520_nn_multiplication: nn_multiplication port map(weight_520 , x_520 ,store_weight_520 );
ut521_nn_multiplication: nn_multiplication port map(weight_521 , x_521 ,store_weight_521 );
ut522_nn_multiplication: nn_multiplication port map(weight_522 , x_522 ,store_weight_522 );
ut523_nn_multiplication: nn_multiplication port map(weight_523 , x_523 ,store_weight_523 );
ut524_nn_multiplication: nn_multiplication port map(weight_524 , x_524 ,store_weight_524 );
ut525_nn_multiplication: nn_multiplication port map(weight_525 , x_525 ,store_weight_525 );
ut526_nn_multiplication: nn_multiplication port map(weight_526 , x_526 ,store_weight_526 );
ut527_nn_multiplication: nn_multiplication port map(weight_527 , x_527 ,store_weight_527 );
ut528_nn_multiplication: nn_multiplication port map(weight_528 , x_528 ,store_weight_528 );
ut529_nn_multiplication: nn_multiplication port map(weight_529 , x_529 ,store_weight_529 );
ut530_nn_multiplication: nn_multiplication port map(weight_530 , x_530 ,store_weight_530 );
ut531_nn_multiplication: nn_multiplication port map(weight_531 , x_531 ,store_weight_531 );
ut532_nn_multiplication: nn_multiplication port map(weight_532 , x_532 ,store_weight_532 );
ut533_nn_multiplication: nn_multiplication port map(weight_533 , x_533 ,store_weight_533 );
ut534_nn_multiplication: nn_multiplication port map(weight_534 , x_534 ,store_weight_534 );
ut535_nn_multiplication: nn_multiplication port map(weight_535 , x_535 ,store_weight_535 );
ut536_nn_multiplication: nn_multiplication port map(weight_536 , x_536 ,store_weight_536 );
ut537_nn_multiplication: nn_multiplication port map(weight_537 , x_537 ,store_weight_537 );
ut538_nn_multiplication: nn_multiplication port map(weight_538 , x_538 ,store_weight_538 );
ut539_nn_multiplication: nn_multiplication port map(weight_539 , x_539 ,store_weight_539 );
ut540_nn_multiplication: nn_multiplication port map(weight_540 , x_540 ,store_weight_540 );
ut541_nn_multiplication: nn_multiplication port map(weight_541 , x_541 ,store_weight_541 );
ut542_nn_multiplication: nn_multiplication port map(weight_542 , x_542 ,store_weight_542 );
ut543_nn_multiplication: nn_multiplication port map(weight_543 , x_543 ,store_weight_543 );
ut544_nn_multiplication: nn_multiplication port map(weight_544 , x_544 ,store_weight_544 );
ut545_nn_multiplication: nn_multiplication port map(weight_545 , x_545 ,store_weight_545 );
ut546_nn_multiplication: nn_multiplication port map(weight_546 , x_546 ,store_weight_546 );
ut547_nn_multiplication: nn_multiplication port map(weight_547 , x_547 ,store_weight_547 );
ut548_nn_multiplication: nn_multiplication port map(weight_548 , x_548 ,store_weight_548 );
ut549_nn_multiplication: nn_multiplication port map(weight_549 , x_549 ,store_weight_549 );
ut550_nn_multiplication: nn_multiplication port map(weight_550 , x_550 ,store_weight_550 );
ut551_nn_multiplication: nn_multiplication port map(weight_551 , x_551 ,store_weight_551 );
ut552_nn_multiplication: nn_multiplication port map(weight_552 , x_552 ,store_weight_552 );
ut553_nn_multiplication: nn_multiplication port map(weight_553 , x_553 ,store_weight_553 );
ut554_nn_multiplication: nn_multiplication port map(weight_554 , x_554 ,store_weight_554 );
ut555_nn_multiplication: nn_multiplication port map(weight_555 , x_555 ,store_weight_555 );
ut556_nn_multiplication: nn_multiplication port map(weight_556 , x_556 ,store_weight_556 );
ut557_nn_multiplication: nn_multiplication port map(weight_557 , x_557 ,store_weight_557 );
ut558_nn_multiplication: nn_multiplication port map(weight_558 , x_558 ,store_weight_558 );
ut559_nn_multiplication: nn_multiplication port map(weight_559 , x_559 ,store_weight_559 );
ut560_nn_multiplication: nn_multiplication port map(weight_560 , x_560 ,store_weight_560 );
ut561_nn_multiplication: nn_multiplication port map(weight_561 , x_561 ,store_weight_561 );
ut562_nn_multiplication: nn_multiplication port map(weight_562 , x_562 ,store_weight_562 );
ut563_nn_multiplication: nn_multiplication port map(weight_563 , x_563 ,store_weight_563 );
ut564_nn_multiplication: nn_multiplication port map(weight_564 , x_564 ,store_weight_564 );
ut565_nn_multiplication: nn_multiplication port map(weight_565 , x_565 ,store_weight_565 );
ut566_nn_multiplication: nn_multiplication port map(weight_566 , x_566 ,store_weight_566 );
ut567_nn_multiplication: nn_multiplication port map(weight_567 , x_567 ,store_weight_567 );
ut568_nn_multiplication: nn_multiplication port map(weight_568 , x_568 ,store_weight_568 );
ut569_nn_multiplication: nn_multiplication port map(weight_569 , x_569 ,store_weight_569 );
ut570_nn_multiplication: nn_multiplication port map(weight_570 , x_570 ,store_weight_570 );
ut571_nn_multiplication: nn_multiplication port map(weight_571 , x_571 ,store_weight_571 );
ut572_nn_multiplication: nn_multiplication port map(weight_572 , x_572 ,store_weight_572 );
ut573_nn_multiplication: nn_multiplication port map(weight_573 , x_573 ,store_weight_573 );
ut574_nn_multiplication: nn_multiplication port map(weight_574 , x_574 ,store_weight_574 );
ut575_nn_multiplication: nn_multiplication port map(weight_575 , x_575 ,store_weight_575 );
ut576_nn_multiplication: nn_multiplication port map(weight_576 , x_576 ,store_weight_576 );
ut577_nn_multiplication: nn_multiplication port map(weight_577 , x_577 ,store_weight_577 );
ut578_nn_multiplication: nn_multiplication port map(weight_578 , x_578 ,store_weight_578 );
ut579_nn_multiplication: nn_multiplication port map(weight_579 , x_579 ,store_weight_579 );
ut580_nn_multiplication: nn_multiplication port map(weight_580 , x_580 ,store_weight_580 );
ut581_nn_multiplication: nn_multiplication port map(weight_581 , x_581 ,store_weight_581 );
ut582_nn_multiplication: nn_multiplication port map(weight_582 , x_582 ,store_weight_582 );
ut583_nn_multiplication: nn_multiplication port map(weight_583 , x_583 ,store_weight_583 );
ut584_nn_multiplication: nn_multiplication port map(weight_584 , x_584 ,store_weight_584 );
ut585_nn_multiplication: nn_multiplication port map(weight_585 , x_585 ,store_weight_585 );
ut586_nn_multiplication: nn_multiplication port map(weight_586 , x_586 ,store_weight_586 );
ut587_nn_multiplication: nn_multiplication port map(weight_587 , x_587 ,store_weight_587 );
ut588_nn_multiplication: nn_multiplication port map(weight_588 , x_588 ,store_weight_588 );
ut589_nn_multiplication: nn_multiplication port map(weight_589 , x_589 ,store_weight_589 );
ut590_nn_multiplication: nn_multiplication port map(weight_590 , x_590 ,store_weight_590 );
ut591_nn_multiplication: nn_multiplication port map(weight_591 , x_591 ,store_weight_591 );
ut592_nn_multiplication: nn_multiplication port map(weight_592 , x_592 ,store_weight_592 );
ut593_nn_multiplication: nn_multiplication port map(weight_593 , x_593 ,store_weight_593 );
ut594_nn_multiplication: nn_multiplication port map(weight_594 , x_594 ,store_weight_594 );
ut595_nn_multiplication: nn_multiplication port map(weight_595 , x_595 ,store_weight_595 );
ut596_nn_multiplication: nn_multiplication port map(weight_596 , x_596 ,store_weight_596 );
ut597_nn_multiplication: nn_multiplication port map(weight_597 , x_597 ,store_weight_597 );
ut598_nn_multiplication: nn_multiplication port map(weight_598 , x_598 ,store_weight_598 );
ut599_nn_multiplication: nn_multiplication port map(weight_599 , x_599 ,store_weight_599 );
ut600_nn_multiplication: nn_multiplication port map(weight_600 , x_600 ,store_weight_600 );
ut601_nn_multiplication: nn_multiplication port map(weight_601 , x_601 ,store_weight_601 );
ut602_nn_multiplication: nn_multiplication port map(weight_602 , x_602 ,store_weight_602 );
ut603_nn_multiplication: nn_multiplication port map(weight_603 , x_603 ,store_weight_603 );
ut604_nn_multiplication: nn_multiplication port map(weight_604 , x_604 ,store_weight_604 );
ut605_nn_multiplication: nn_multiplication port map(weight_605 , x_605 ,store_weight_605 );
ut606_nn_multiplication: nn_multiplication port map(weight_606 , x_606 ,store_weight_606 );
ut607_nn_multiplication: nn_multiplication port map(weight_607 , x_607 ,store_weight_607 );
ut608_nn_multiplication: nn_multiplication port map(weight_608 , x_608 ,store_weight_608 );
ut609_nn_multiplication: nn_multiplication port map(weight_609 , x_609 ,store_weight_609 );
ut610_nn_multiplication: nn_multiplication port map(weight_610 , x_610 ,store_weight_610 );
ut611_nn_multiplication: nn_multiplication port map(weight_611 , x_611 ,store_weight_611 );
ut612_nn_multiplication: nn_multiplication port map(weight_612 , x_612 ,store_weight_612 );
ut613_nn_multiplication: nn_multiplication port map(weight_613 , x_613 ,store_weight_613 );
ut614_nn_multiplication: nn_multiplication port map(weight_614 , x_614 ,store_weight_614 );
ut615_nn_multiplication: nn_multiplication port map(weight_615 , x_615 ,store_weight_615 );
ut616_nn_multiplication: nn_multiplication port map(weight_616 , x_616 ,store_weight_616 );
ut617_nn_multiplication: nn_multiplication port map(weight_617 , x_617 ,store_weight_617 );
ut618_nn_multiplication: nn_multiplication port map(weight_618 , x_618 ,store_weight_618 );
ut619_nn_multiplication: nn_multiplication port map(weight_619 , x_619 ,store_weight_619 );
ut620_nn_multiplication: nn_multiplication port map(weight_620 , x_620 ,store_weight_620 );
ut621_nn_multiplication: nn_multiplication port map(weight_621 , x_621 ,store_weight_621 );
ut622_nn_multiplication: nn_multiplication port map(weight_622 , x_622 ,store_weight_622 );
ut623_nn_multiplication: nn_multiplication port map(weight_623 , x_623 ,store_weight_623 );
ut624_nn_multiplication: nn_multiplication port map(weight_624 , x_624 ,store_weight_624 );
ut625_nn_multiplication: nn_multiplication port map(weight_625 , x_625 ,store_weight_625 );
ut626_nn_multiplication: nn_multiplication port map(weight_626 , x_626 ,store_weight_626 );
ut627_nn_multiplication: nn_multiplication port map(weight_627 , x_627 ,store_weight_627 );
ut628_nn_multiplication: nn_multiplication port map(weight_628 , x_628 ,store_weight_628 );
ut629_nn_multiplication: nn_multiplication port map(weight_629 , x_629 ,store_weight_629 );
ut630_nn_multiplication: nn_multiplication port map(weight_630 , x_630 ,store_weight_630 );
ut631_nn_multiplication: nn_multiplication port map(weight_631 , x_631 ,store_weight_631 );
ut632_nn_multiplication: nn_multiplication port map(weight_632 , x_632 ,store_weight_632 );
ut633_nn_multiplication: nn_multiplication port map(weight_633 , x_633 ,store_weight_633 );
ut634_nn_multiplication: nn_multiplication port map(weight_634 , x_634 ,store_weight_634 );
ut635_nn_multiplication: nn_multiplication port map(weight_635 , x_635 ,store_weight_635 );
ut636_nn_multiplication: nn_multiplication port map(weight_636 , x_636 ,store_weight_636 );
ut637_nn_multiplication: nn_multiplication port map(weight_637 , x_637 ,store_weight_637 );
ut638_nn_multiplication: nn_multiplication port map(weight_638 , x_638 ,store_weight_638 );
ut639_nn_multiplication: nn_multiplication port map(weight_639 , x_639 ,store_weight_639 );
ut640_nn_multiplication: nn_multiplication port map(weight_640 , x_640 ,store_weight_640 );
ut641_nn_multiplication: nn_multiplication port map(weight_641 , x_641 ,store_weight_641 );
ut642_nn_multiplication: nn_multiplication port map(weight_642 , x_642 ,store_weight_642 );
ut643_nn_multiplication: nn_multiplication port map(weight_643 , x_643 ,store_weight_643 );
ut644_nn_multiplication: nn_multiplication port map(weight_644 , x_644 ,store_weight_644 );
ut645_nn_multiplication: nn_multiplication port map(weight_645 , x_645 ,store_weight_645 );
ut646_nn_multiplication: nn_multiplication port map(weight_646 , x_646 ,store_weight_646 );
ut647_nn_multiplication: nn_multiplication port map(weight_647 , x_647 ,store_weight_647 );
ut648_nn_multiplication: nn_multiplication port map(weight_648 , x_648 ,store_weight_648 );
ut649_nn_multiplication: nn_multiplication port map(weight_649 , x_649 ,store_weight_649 );
ut650_nn_multiplication: nn_multiplication port map(weight_650 , x_650 ,store_weight_650 );
ut651_nn_multiplication: nn_multiplication port map(weight_651 , x_651 ,store_weight_651 );
ut652_nn_multiplication: nn_multiplication port map(weight_652 , x_652 ,store_weight_652 );
ut653_nn_multiplication: nn_multiplication port map(weight_653 , x_653 ,store_weight_653 );
ut654_nn_multiplication: nn_multiplication port map(weight_654 , x_654 ,store_weight_654 );
ut655_nn_multiplication: nn_multiplication port map(weight_655 , x_655 ,store_weight_655 );
ut656_nn_multiplication: nn_multiplication port map(weight_656 , x_656 ,store_weight_656 );
ut657_nn_multiplication: nn_multiplication port map(weight_657 , x_657 ,store_weight_657 );
ut658_nn_multiplication: nn_multiplication port map(weight_658 , x_658 ,store_weight_658 );
ut659_nn_multiplication: nn_multiplication port map(weight_659 , x_659 ,store_weight_659 );
ut660_nn_multiplication: nn_multiplication port map(weight_660 , x_660 ,store_weight_660 );
ut661_nn_multiplication: nn_multiplication port map(weight_661 , x_661 ,store_weight_661 );
ut662_nn_multiplication: nn_multiplication port map(weight_662 , x_662 ,store_weight_662 );
ut663_nn_multiplication: nn_multiplication port map(weight_663 , x_663 ,store_weight_663 );
ut664_nn_multiplication: nn_multiplication port map(weight_664 , x_664 ,store_weight_664 );
ut665_nn_multiplication: nn_multiplication port map(weight_665 , x_665 ,store_weight_665 );
ut666_nn_multiplication: nn_multiplication port map(weight_666 , x_666 ,store_weight_666 );
ut667_nn_multiplication: nn_multiplication port map(weight_667 , x_667 ,store_weight_667 );
ut668_nn_multiplication: nn_multiplication port map(weight_668 , x_668 ,store_weight_668 );
ut669_nn_multiplication: nn_multiplication port map(weight_669 , x_669 ,store_weight_669 );
ut670_nn_multiplication: nn_multiplication port map(weight_670 , x_670 ,store_weight_670 );
ut671_nn_multiplication: nn_multiplication port map(weight_671 , x_671 ,store_weight_671 );
ut672_nn_multiplication: nn_multiplication port map(weight_672 , x_672 ,store_weight_672 );
ut673_nn_multiplication: nn_multiplication port map(weight_673 , x_673 ,store_weight_673 );
ut674_nn_multiplication: nn_multiplication port map(weight_674 , x_674 ,store_weight_674 );
ut675_nn_multiplication: nn_multiplication port map(weight_675 , x_675 ,store_weight_675 );
ut676_nn_multiplication: nn_multiplication port map(weight_676 , x_676 ,store_weight_676 );
ut677_nn_multiplication: nn_multiplication port map(weight_677 , x_677 ,store_weight_677 );
ut678_nn_multiplication: nn_multiplication port map(weight_678 , x_678 ,store_weight_678 );
ut679_nn_multiplication: nn_multiplication port map(weight_679 , x_679 ,store_weight_679 );
ut680_nn_multiplication: nn_multiplication port map(weight_680 , x_680 ,store_weight_680 );
ut681_nn_multiplication: nn_multiplication port map(weight_681 , x_681 ,store_weight_681 );
ut682_nn_multiplication: nn_multiplication port map(weight_682 , x_682 ,store_weight_682 );
ut683_nn_multiplication: nn_multiplication port map(weight_683 , x_683 ,store_weight_683 );
ut684_nn_multiplication: nn_multiplication port map(weight_684 , x_684 ,store_weight_684 );
ut685_nn_multiplication: nn_multiplication port map(weight_685 , x_685 ,store_weight_685 );
ut686_nn_multiplication: nn_multiplication port map(weight_686 , x_686 ,store_weight_686 );
ut687_nn_multiplication: nn_multiplication port map(weight_687 , x_687 ,store_weight_687 );
ut688_nn_multiplication: nn_multiplication port map(weight_688 , x_688 ,store_weight_688 );
ut689_nn_multiplication: nn_multiplication port map(weight_689 , x_689 ,store_weight_689 );
ut690_nn_multiplication: nn_multiplication port map(weight_690 , x_690 ,store_weight_690 );
ut691_nn_multiplication: nn_multiplication port map(weight_691 , x_691 ,store_weight_691 );
ut692_nn_multiplication: nn_multiplication port map(weight_692 , x_692 ,store_weight_692 );
ut693_nn_multiplication: nn_multiplication port map(weight_693 , x_693 ,store_weight_693 );
ut694_nn_multiplication: nn_multiplication port map(weight_694 , x_694 ,store_weight_694 );
ut695_nn_multiplication: nn_multiplication port map(weight_695 , x_695 ,store_weight_695 );
ut696_nn_multiplication: nn_multiplication port map(weight_696 , x_696 ,store_weight_696 );
ut697_nn_multiplication: nn_multiplication port map(weight_697 , x_697 ,store_weight_697 );
ut698_nn_multiplication: nn_multiplication port map(weight_698 , x_698 ,store_weight_698 );
ut699_nn_multiplication: nn_multiplication port map(weight_699 , x_699 ,store_weight_699 );
ut700_nn_multiplication: nn_multiplication port map(weight_700 , x_700 ,store_weight_700 );
ut701_nn_multiplication: nn_multiplication port map(weight_701 , x_701 ,store_weight_701 );
ut702_nn_multiplication: nn_multiplication port map(weight_702 , x_702 ,store_weight_702 );
ut703_nn_multiplication: nn_multiplication port map(weight_703 , x_703 ,store_weight_703 );
ut704_nn_multiplication: nn_multiplication port map(weight_704 , x_704 ,store_weight_704 );
ut705_nn_multiplication: nn_multiplication port map(weight_705 , x_705 ,store_weight_705 );
ut706_nn_multiplication: nn_multiplication port map(weight_706 , x_706 ,store_weight_706 );
ut707_nn_multiplication: nn_multiplication port map(weight_707 , x_707 ,store_weight_707 );
ut708_nn_multiplication: nn_multiplication port map(weight_708 , x_708 ,store_weight_708 );
ut709_nn_multiplication: nn_multiplication port map(weight_709 , x_709 ,store_weight_709 );
ut710_nn_multiplication: nn_multiplication port map(weight_710 , x_710 ,store_weight_710 );
ut711_nn_multiplication: nn_multiplication port map(weight_711 , x_711 ,store_weight_711 );
ut712_nn_multiplication: nn_multiplication port map(weight_712 , x_712 ,store_weight_712 );
ut713_nn_multiplication: nn_multiplication port map(weight_713 , x_713 ,store_weight_713 );
ut714_nn_multiplication: nn_multiplication port map(weight_714 , x_714 ,store_weight_714 );
ut715_nn_multiplication: nn_multiplication port map(weight_715 , x_715 ,store_weight_715 );
ut716_nn_multiplication: nn_multiplication port map(weight_716 , x_716 ,store_weight_716 );
ut717_nn_multiplication: nn_multiplication port map(weight_717 , x_717 ,store_weight_717 );
ut718_nn_multiplication: nn_multiplication port map(weight_718 , x_718 ,store_weight_718 );
ut719_nn_multiplication: nn_multiplication port map(weight_719 , x_719 ,store_weight_719 );
ut720_nn_multiplication: nn_multiplication port map(weight_720 , x_720 ,store_weight_720 );
ut721_nn_multiplication: nn_multiplication port map(weight_721 , x_721 ,store_weight_721 );
ut722_nn_multiplication: nn_multiplication port map(weight_722 , x_722 ,store_weight_722 );
ut723_nn_multiplication: nn_multiplication port map(weight_723 , x_723 ,store_weight_723 );
ut724_nn_multiplication: nn_multiplication port map(weight_724 , x_724 ,store_weight_724 );
ut725_nn_multiplication: nn_multiplication port map(weight_725 , x_725 ,store_weight_725 );
ut726_nn_multiplication: nn_multiplication port map(weight_726 , x_726 ,store_weight_726 );
ut727_nn_multiplication: nn_multiplication port map(weight_727 , x_727 ,store_weight_727 );
ut728_nn_multiplication: nn_multiplication port map(weight_728 , x_728 ,store_weight_728 );
ut729_nn_multiplication: nn_multiplication port map(weight_729 , x_729 ,store_weight_729 );
ut730_nn_multiplication: nn_multiplication port map(weight_730 , x_730 ,store_weight_730 );
ut731_nn_multiplication: nn_multiplication port map(weight_731 , x_731 ,store_weight_731 );
ut732_nn_multiplication: nn_multiplication port map(weight_732 , x_732 ,store_weight_732 );
ut733_nn_multiplication: nn_multiplication port map(weight_733 , x_733 ,store_weight_733 );
ut734_nn_multiplication: nn_multiplication port map(weight_734 , x_734 ,store_weight_734 );
ut735_nn_multiplication: nn_multiplication port map(weight_735 , x_735 ,store_weight_735 );
ut736_nn_multiplication: nn_multiplication port map(weight_736 , x_736 ,store_weight_736 );
ut737_nn_multiplication: nn_multiplication port map(weight_737 , x_737 ,store_weight_737 );
ut738_nn_multiplication: nn_multiplication port map(weight_738 , x_738 ,store_weight_738 );
ut739_nn_multiplication: nn_multiplication port map(weight_739 , x_739 ,store_weight_739 );
ut740_nn_multiplication: nn_multiplication port map(weight_740 , x_740 ,store_weight_740 );
ut741_nn_multiplication: nn_multiplication port map(weight_741 , x_741 ,store_weight_741 );
ut742_nn_multiplication: nn_multiplication port map(weight_742 , x_742 ,store_weight_742 );
ut743_nn_multiplication: nn_multiplication port map(weight_743 , x_743 ,store_weight_743 );
ut744_nn_multiplication: nn_multiplication port map(weight_744 , x_744 ,store_weight_744 );
ut745_nn_multiplication: nn_multiplication port map(weight_745 , x_745 ,store_weight_745 );
ut746_nn_multiplication: nn_multiplication port map(weight_746 , x_746 ,store_weight_746 );
ut747_nn_multiplication: nn_multiplication port map(weight_747 , x_747 ,store_weight_747 );
ut748_nn_multiplication: nn_multiplication port map(weight_748 , x_748 ,store_weight_748 );
ut749_nn_multiplication: nn_multiplication port map(weight_749 , x_749 ,store_weight_749 );
ut750_nn_multiplication: nn_multiplication port map(weight_750 , x_750 ,store_weight_750 );
ut751_nn_multiplication: nn_multiplication port map(weight_751 , x_751 ,store_weight_751 );
ut752_nn_multiplication: nn_multiplication port map(weight_752 , x_752 ,store_weight_752 );
ut753_nn_multiplication: nn_multiplication port map(weight_753 , x_753 ,store_weight_753 );
ut754_nn_multiplication: nn_multiplication port map(weight_754 , x_754 ,store_weight_754 );
ut755_nn_multiplication: nn_multiplication port map(weight_755 , x_755 ,store_weight_755 );
ut756_nn_multiplication: nn_multiplication port map(weight_756 , x_756 ,store_weight_756 );
ut757_nn_multiplication: nn_multiplication port map(weight_757 , x_757 ,store_weight_757 );
ut758_nn_multiplication: nn_multiplication port map(weight_758 , x_758 ,store_weight_758 );
ut759_nn_multiplication: nn_multiplication port map(weight_759 , x_759 ,store_weight_759 );
ut760_nn_multiplication: nn_multiplication port map(weight_760 , x_760 ,store_weight_760 );
ut761_nn_multiplication: nn_multiplication port map(weight_761 , x_761 ,store_weight_761 );
ut762_nn_multiplication: nn_multiplication port map(weight_762 , x_762 ,store_weight_762 );
ut763_nn_multiplication: nn_multiplication port map(weight_763 , x_763 ,store_weight_763 );
ut764_nn_multiplication: nn_multiplication port map(weight_764 , x_764 ,store_weight_764 );
ut765_nn_multiplication: nn_multiplication port map(weight_765 , x_765 ,store_weight_765 );
ut766_nn_multiplication: nn_multiplication port map(weight_766 , x_766 ,store_weight_766 );
ut767_nn_multiplication: nn_multiplication port map(weight_767 , x_767 ,store_weight_767 );
ut768_nn_multiplication: nn_multiplication port map(weight_768 , x_768 ,store_weight_768 );
ut769_nn_multiplication: nn_multiplication port map(weight_769 , x_769 ,store_weight_769 );
ut770_nn_multiplication: nn_multiplication port map(weight_770 , x_770 ,store_weight_770 );
ut771_nn_multiplication: nn_multiplication port map(weight_771 , x_771 ,store_weight_771 );
ut772_nn_multiplication: nn_multiplication port map(weight_772 , x_772 ,store_weight_772 );
ut773_nn_multiplication: nn_multiplication port map(weight_773 , x_773 ,store_weight_773 );
ut774_nn_multiplication: nn_multiplication port map(weight_774 , x_774 ,store_weight_774 );
ut775_nn_multiplication: nn_multiplication port map(weight_775 , x_775 ,store_weight_775 );
ut776_nn_multiplication: nn_multiplication port map(weight_776 , x_776 ,store_weight_776 );
ut777_nn_multiplication: nn_multiplication port map(weight_777 , x_777 ,store_weight_777 );
ut778_nn_multiplication: nn_multiplication port map(weight_778 , x_778 ,store_weight_778 );
ut779_nn_multiplication: nn_multiplication port map(weight_779 , x_779 ,store_weight_779 );
ut780_nn_multiplication: nn_multiplication port map(weight_780 , x_780 ,store_weight_780 );
ut781_nn_multiplication: nn_multiplication port map(weight_781 , x_781 ,store_weight_781 );
ut782_nn_multiplication: nn_multiplication port map(weight_782 , x_782 ,store_weight_782 );
ut783_nn_multiplication: nn_multiplication port map(weight_783 , x_783 ,store_weight_783 );
ut0_nn_addition: nn_addition port map( store_weight_0,store_weight_1,sum_0);
ut1_nn_addition: nn_addition port map( store_weight_2,store_weight_3,sum_1);
ut2_nn_addition: nn_addition port map( store_weight_4,store_weight_5,sum_2);
ut3_nn_addition: nn_addition port map( store_weight_6,store_weight_7,sum_3);
ut4_nn_addition: nn_addition port map( store_weight_8,store_weight_9,sum_4);
ut5_nn_addition: nn_addition port map( store_weight_10,store_weight_11,sum_5);
ut6_nn_addition: nn_addition port map( store_weight_12,store_weight_13,sum_6);
ut7_nn_addition: nn_addition port map( store_weight_14,store_weight_15,sum_7);
ut8_nn_addition: nn_addition port map( store_weight_16,store_weight_17,sum_8);
ut9_nn_addition: nn_addition port map( store_weight_18,store_weight_19,sum_9);
ut10_nn_addition: nn_addition port map( store_weight_20,store_weight_21,sum_10);
ut11_nn_addition: nn_addition port map( store_weight_22,store_weight_23,sum_11);
ut12_nn_addition: nn_addition port map( store_weight_24,store_weight_25,sum_12);
ut13_nn_addition: nn_addition port map( store_weight_26,store_weight_27,sum_13);
ut14_nn_addition: nn_addition port map( store_weight_28,store_weight_29,sum_14);
ut15_nn_addition: nn_addition port map( store_weight_30,store_weight_31,sum_15);
ut16_nn_addition: nn_addition port map( store_weight_32,store_weight_33,sum_16);
ut17_nn_addition: nn_addition port map( store_weight_34,store_weight_35,sum_17);
ut18_nn_addition: nn_addition port map( store_weight_36,store_weight_37,sum_18);
ut19_nn_addition: nn_addition port map( store_weight_38,store_weight_39,sum_19);
ut20_nn_addition: nn_addition port map( store_weight_40,store_weight_41,sum_20);
ut21_nn_addition: nn_addition port map( store_weight_42,store_weight_43,sum_21);
ut22_nn_addition: nn_addition port map( store_weight_44,store_weight_45,sum_22);
ut23_nn_addition: nn_addition port map( store_weight_46,store_weight_47,sum_23);
ut24_nn_addition: nn_addition port map( store_weight_48,store_weight_49,sum_24);
ut25_nn_addition: nn_addition port map( store_weight_50,store_weight_51,sum_25);
ut26_nn_addition: nn_addition port map( store_weight_52,store_weight_53,sum_26);
ut27_nn_addition: nn_addition port map( store_weight_54,store_weight_55,sum_27);
ut28_nn_addition: nn_addition port map( store_weight_56,store_weight_57,sum_28);
ut29_nn_addition: nn_addition port map( store_weight_58,store_weight_59,sum_29);
ut30_nn_addition: nn_addition port map( store_weight_60,store_weight_61,sum_30);
ut31_nn_addition: nn_addition port map( store_weight_62,store_weight_63,sum_31);
ut32_nn_addition: nn_addition port map( store_weight_64,store_weight_65,sum_32);
ut33_nn_addition: nn_addition port map( store_weight_66,store_weight_67,sum_33);
ut34_nn_addition: nn_addition port map( store_weight_68,store_weight_69,sum_34);
ut35_nn_addition: nn_addition port map( store_weight_70,store_weight_71,sum_35);
ut36_nn_addition: nn_addition port map( store_weight_72,store_weight_73,sum_36);
ut37_nn_addition: nn_addition port map( store_weight_74,store_weight_75,sum_37);
ut38_nn_addition: nn_addition port map( store_weight_76,store_weight_77,sum_38);
ut39_nn_addition: nn_addition port map( store_weight_78,store_weight_79,sum_39);
ut40_nn_addition: nn_addition port map( store_weight_80,store_weight_81,sum_40);
ut41_nn_addition: nn_addition port map( store_weight_82,store_weight_83,sum_41);
ut42_nn_addition: nn_addition port map( store_weight_84,store_weight_85,sum_42);
ut43_nn_addition: nn_addition port map( store_weight_86,store_weight_87,sum_43);
ut44_nn_addition: nn_addition port map( store_weight_88,store_weight_89,sum_44);
ut45_nn_addition: nn_addition port map( store_weight_90,store_weight_91,sum_45);
ut46_nn_addition: nn_addition port map( store_weight_92,store_weight_93,sum_46);
ut47_nn_addition: nn_addition port map( store_weight_94,store_weight_95,sum_47);
ut48_nn_addition: nn_addition port map( store_weight_96,store_weight_97,sum_48);
ut49_nn_addition: nn_addition port map( store_weight_98,store_weight_99,sum_49);
ut50_nn_addition: nn_addition port map( store_weight_100,store_weight_101,sum_50);
ut51_nn_addition: nn_addition port map( store_weight_102,store_weight_103,sum_51);
ut52_nn_addition: nn_addition port map( store_weight_104,store_weight_105,sum_52);
ut53_nn_addition: nn_addition port map( store_weight_106,store_weight_107,sum_53);
ut54_nn_addition: nn_addition port map( store_weight_108,store_weight_109,sum_54);
ut55_nn_addition: nn_addition port map( store_weight_110,store_weight_111,sum_55);
ut56_nn_addition: nn_addition port map( store_weight_112,store_weight_113,sum_56);
ut57_nn_addition: nn_addition port map( store_weight_114,store_weight_115,sum_57);
ut58_nn_addition: nn_addition port map( store_weight_116,store_weight_117,sum_58);
ut59_nn_addition: nn_addition port map( store_weight_118,store_weight_119,sum_59);
ut60_nn_addition: nn_addition port map( store_weight_120,store_weight_121,sum_60);
ut61_nn_addition: nn_addition port map( store_weight_122,store_weight_123,sum_61);
ut62_nn_addition: nn_addition port map( store_weight_124,store_weight_125,sum_62);
ut63_nn_addition: nn_addition port map( store_weight_126,store_weight_127,sum_63);
ut64_nn_addition: nn_addition port map( store_weight_128,store_weight_129,sum_64);
ut65_nn_addition: nn_addition port map( store_weight_130,store_weight_131,sum_65);
ut66_nn_addition: nn_addition port map( store_weight_132,store_weight_133,sum_66);
ut67_nn_addition: nn_addition port map( store_weight_134,store_weight_135,sum_67);
ut68_nn_addition: nn_addition port map( store_weight_136,store_weight_137,sum_68);
ut69_nn_addition: nn_addition port map( store_weight_138,store_weight_139,sum_69);
ut70_nn_addition: nn_addition port map( store_weight_140,store_weight_141,sum_70);
ut71_nn_addition: nn_addition port map( store_weight_142,store_weight_143,sum_71);
ut72_nn_addition: nn_addition port map( store_weight_144,store_weight_145,sum_72);
ut73_nn_addition: nn_addition port map( store_weight_146,store_weight_147,sum_73);
ut74_nn_addition: nn_addition port map( store_weight_148,store_weight_149,sum_74);
ut75_nn_addition: nn_addition port map( store_weight_150,store_weight_151,sum_75);
ut76_nn_addition: nn_addition port map( store_weight_152,store_weight_153,sum_76);
ut77_nn_addition: nn_addition port map( store_weight_154,store_weight_155,sum_77);
ut78_nn_addition: nn_addition port map( store_weight_156,store_weight_157,sum_78);
ut79_nn_addition: nn_addition port map( store_weight_158,store_weight_159,sum_79);
ut80_nn_addition: nn_addition port map( store_weight_160,store_weight_161,sum_80);
ut81_nn_addition: nn_addition port map( store_weight_162,store_weight_163,sum_81);
ut82_nn_addition: nn_addition port map( store_weight_164,store_weight_165,sum_82);
ut83_nn_addition: nn_addition port map( store_weight_166,store_weight_167,sum_83);
ut84_nn_addition: nn_addition port map( store_weight_168,store_weight_169,sum_84);
ut85_nn_addition: nn_addition port map( store_weight_170,store_weight_171,sum_85);
ut86_nn_addition: nn_addition port map( store_weight_172,store_weight_173,sum_86);
ut87_nn_addition: nn_addition port map( store_weight_174,store_weight_175,sum_87);
ut88_nn_addition: nn_addition port map( store_weight_176,store_weight_177,sum_88);
ut89_nn_addition: nn_addition port map( store_weight_178,store_weight_179,sum_89);
ut90_nn_addition: nn_addition port map( store_weight_180,store_weight_181,sum_90);
ut91_nn_addition: nn_addition port map( store_weight_182,store_weight_183,sum_91);
ut92_nn_addition: nn_addition port map( store_weight_184,store_weight_185,sum_92);
ut93_nn_addition: nn_addition port map( store_weight_186,store_weight_187,sum_93);
ut94_nn_addition: nn_addition port map( store_weight_188,store_weight_189,sum_94);
ut95_nn_addition: nn_addition port map( store_weight_190,store_weight_191,sum_95);
ut96_nn_addition: nn_addition port map( store_weight_192,store_weight_193,sum_96);
ut97_nn_addition: nn_addition port map( store_weight_194,store_weight_195,sum_97);
ut98_nn_addition: nn_addition port map( store_weight_196,store_weight_197,sum_98);
ut99_nn_addition: nn_addition port map( store_weight_198,store_weight_199,sum_99);
ut100_nn_addition: nn_addition port map( store_weight_200,store_weight_201,sum_100);
ut101_nn_addition: nn_addition port map( store_weight_202,store_weight_203,sum_101);
ut102_nn_addition: nn_addition port map( store_weight_204,store_weight_205,sum_102);
ut103_nn_addition: nn_addition port map( store_weight_206,store_weight_207,sum_103);
ut104_nn_addition: nn_addition port map( store_weight_208,store_weight_209,sum_104);
ut105_nn_addition: nn_addition port map( store_weight_210,store_weight_211,sum_105);
ut106_nn_addition: nn_addition port map( store_weight_212,store_weight_213,sum_106);
ut107_nn_addition: nn_addition port map( store_weight_214,store_weight_215,sum_107);
ut108_nn_addition: nn_addition port map( store_weight_216,store_weight_217,sum_108);
ut109_nn_addition: nn_addition port map( store_weight_218,store_weight_219,sum_109);
ut110_nn_addition: nn_addition port map( store_weight_220,store_weight_221,sum_110);
ut111_nn_addition: nn_addition port map( store_weight_222,store_weight_223,sum_111);
ut112_nn_addition: nn_addition port map( store_weight_224,store_weight_225,sum_112);
ut113_nn_addition: nn_addition port map( store_weight_226,store_weight_227,sum_113);
ut114_nn_addition: nn_addition port map( store_weight_228,store_weight_229,sum_114);
ut115_nn_addition: nn_addition port map( store_weight_230,store_weight_231,sum_115);
ut116_nn_addition: nn_addition port map( store_weight_232,store_weight_233,sum_116);
ut117_nn_addition: nn_addition port map( store_weight_234,store_weight_235,sum_117);
ut118_nn_addition: nn_addition port map( store_weight_236,store_weight_237,sum_118);
ut119_nn_addition: nn_addition port map( store_weight_238,store_weight_239,sum_119);
ut120_nn_addition: nn_addition port map( store_weight_240,store_weight_241,sum_120);
ut121_nn_addition: nn_addition port map( store_weight_242,store_weight_243,sum_121);
ut122_nn_addition: nn_addition port map( store_weight_244,store_weight_245,sum_122);
ut123_nn_addition: nn_addition port map( store_weight_246,store_weight_247,sum_123);
ut124_nn_addition: nn_addition port map( store_weight_248,store_weight_249,sum_124);
ut125_nn_addition: nn_addition port map( store_weight_250,store_weight_251,sum_125);
ut126_nn_addition: nn_addition port map( store_weight_252,store_weight_253,sum_126);
ut127_nn_addition: nn_addition port map( store_weight_254,store_weight_255,sum_127);
ut128_nn_addition: nn_addition port map( store_weight_256,store_weight_257,sum_128);
ut129_nn_addition: nn_addition port map( store_weight_258,store_weight_259,sum_129);
ut130_nn_addition: nn_addition port map( store_weight_260,store_weight_261,sum_130);
ut131_nn_addition: nn_addition port map( store_weight_262,store_weight_263,sum_131);
ut132_nn_addition: nn_addition port map( store_weight_264,store_weight_265,sum_132);
ut133_nn_addition: nn_addition port map( store_weight_266,store_weight_267,sum_133);
ut134_nn_addition: nn_addition port map( store_weight_268,store_weight_269,sum_134);
ut135_nn_addition: nn_addition port map( store_weight_270,store_weight_271,sum_135);
ut136_nn_addition: nn_addition port map( store_weight_272,store_weight_273,sum_136);
ut137_nn_addition: nn_addition port map( store_weight_274,store_weight_275,sum_137);
ut138_nn_addition: nn_addition port map( store_weight_276,store_weight_277,sum_138);
ut139_nn_addition: nn_addition port map( store_weight_278,store_weight_279,sum_139);
ut140_nn_addition: nn_addition port map( store_weight_280,store_weight_281,sum_140);
ut141_nn_addition: nn_addition port map( store_weight_282,store_weight_283,sum_141);
ut142_nn_addition: nn_addition port map( store_weight_284,store_weight_285,sum_142);
ut143_nn_addition: nn_addition port map( store_weight_286,store_weight_287,sum_143);
ut144_nn_addition: nn_addition port map( store_weight_288,store_weight_289,sum_144);
ut145_nn_addition: nn_addition port map( store_weight_290,store_weight_291,sum_145);
ut146_nn_addition: nn_addition port map( store_weight_292,store_weight_293,sum_146);
ut147_nn_addition: nn_addition port map( store_weight_294,store_weight_295,sum_147);
ut148_nn_addition: nn_addition port map( store_weight_296,store_weight_297,sum_148);
ut149_nn_addition: nn_addition port map( store_weight_298,store_weight_299,sum_149);
ut150_nn_addition: nn_addition port map( store_weight_300,store_weight_301,sum_150);
ut151_nn_addition: nn_addition port map( store_weight_302,store_weight_303,sum_151);
ut152_nn_addition: nn_addition port map( store_weight_304,store_weight_305,sum_152);
ut153_nn_addition: nn_addition port map( store_weight_306,store_weight_307,sum_153);
ut154_nn_addition: nn_addition port map( store_weight_308,store_weight_309,sum_154);
ut155_nn_addition: nn_addition port map( store_weight_310,store_weight_311,sum_155);
ut156_nn_addition: nn_addition port map( store_weight_312,store_weight_313,sum_156);
ut157_nn_addition: nn_addition port map( store_weight_314,store_weight_315,sum_157);
ut158_nn_addition: nn_addition port map( store_weight_316,store_weight_317,sum_158);
ut159_nn_addition: nn_addition port map( store_weight_318,store_weight_319,sum_159);
ut160_nn_addition: nn_addition port map( store_weight_320,store_weight_321,sum_160);
ut161_nn_addition: nn_addition port map( store_weight_322,store_weight_323,sum_161);
ut162_nn_addition: nn_addition port map( store_weight_324,store_weight_325,sum_162);
ut163_nn_addition: nn_addition port map( store_weight_326,store_weight_327,sum_163);
ut164_nn_addition: nn_addition port map( store_weight_328,store_weight_329,sum_164);
ut165_nn_addition: nn_addition port map( store_weight_330,store_weight_331,sum_165);
ut166_nn_addition: nn_addition port map( store_weight_332,store_weight_333,sum_166);
ut167_nn_addition: nn_addition port map( store_weight_334,store_weight_335,sum_167);
ut168_nn_addition: nn_addition port map( store_weight_336,store_weight_337,sum_168);
ut169_nn_addition: nn_addition port map( store_weight_338,store_weight_339,sum_169);
ut170_nn_addition: nn_addition port map( store_weight_340,store_weight_341,sum_170);
ut171_nn_addition: nn_addition port map( store_weight_342,store_weight_343,sum_171);
ut172_nn_addition: nn_addition port map( store_weight_344,store_weight_345,sum_172);
ut173_nn_addition: nn_addition port map( store_weight_346,store_weight_347,sum_173);
ut174_nn_addition: nn_addition port map( store_weight_348,store_weight_349,sum_174);
ut175_nn_addition: nn_addition port map( store_weight_350,store_weight_351,sum_175);
ut176_nn_addition: nn_addition port map( store_weight_352,store_weight_353,sum_176);
ut177_nn_addition: nn_addition port map( store_weight_354,store_weight_355,sum_177);
ut178_nn_addition: nn_addition port map( store_weight_356,store_weight_357,sum_178);
ut179_nn_addition: nn_addition port map( store_weight_358,store_weight_359,sum_179);
ut180_nn_addition: nn_addition port map( store_weight_360,store_weight_361,sum_180);
ut181_nn_addition: nn_addition port map( store_weight_362,store_weight_363,sum_181);
ut182_nn_addition: nn_addition port map( store_weight_364,store_weight_365,sum_182);
ut183_nn_addition: nn_addition port map( store_weight_366,store_weight_367,sum_183);
ut184_nn_addition: nn_addition port map( store_weight_368,store_weight_369,sum_184);
ut185_nn_addition: nn_addition port map( store_weight_370,store_weight_371,sum_185);
ut186_nn_addition: nn_addition port map( store_weight_372,store_weight_373,sum_186);
ut187_nn_addition: nn_addition port map( store_weight_374,store_weight_375,sum_187);
ut188_nn_addition: nn_addition port map( store_weight_376,store_weight_377,sum_188);
ut189_nn_addition: nn_addition port map( store_weight_378,store_weight_379,sum_189);
ut190_nn_addition: nn_addition port map( store_weight_380,store_weight_381,sum_190);
ut191_nn_addition: nn_addition port map( store_weight_382,store_weight_383,sum_191);
ut192_nn_addition: nn_addition port map( store_weight_384,store_weight_385,sum_192);
ut193_nn_addition: nn_addition port map( store_weight_386,store_weight_387,sum_193);
ut194_nn_addition: nn_addition port map( store_weight_388,store_weight_389,sum_194);
ut195_nn_addition: nn_addition port map( store_weight_390,store_weight_391,sum_195);
ut196_nn_addition: nn_addition port map( store_weight_392,store_weight_393,sum_196);
ut197_nn_addition: nn_addition port map( store_weight_394,store_weight_395,sum_197);
ut198_nn_addition: nn_addition port map( store_weight_396,store_weight_397,sum_198);
ut199_nn_addition: nn_addition port map( store_weight_398,store_weight_399,sum_199);
ut200_nn_addition: nn_addition port map( store_weight_400,store_weight_401,sum_200);
ut201_nn_addition: nn_addition port map( store_weight_402,store_weight_403,sum_201);
ut202_nn_addition: nn_addition port map( store_weight_404,store_weight_405,sum_202);
ut203_nn_addition: nn_addition port map( store_weight_406,store_weight_407,sum_203);
ut204_nn_addition: nn_addition port map( store_weight_408,store_weight_409,sum_204);
ut205_nn_addition: nn_addition port map( store_weight_410,store_weight_411,sum_205);
ut206_nn_addition: nn_addition port map( store_weight_412,store_weight_413,sum_206);
ut207_nn_addition: nn_addition port map( store_weight_414,store_weight_415,sum_207);
ut208_nn_addition: nn_addition port map( store_weight_416,store_weight_417,sum_208);
ut209_nn_addition: nn_addition port map( store_weight_418,store_weight_419,sum_209);
ut210_nn_addition: nn_addition port map( store_weight_420,store_weight_421,sum_210);
ut211_nn_addition: nn_addition port map( store_weight_422,store_weight_423,sum_211);
ut212_nn_addition: nn_addition port map( store_weight_424,store_weight_425,sum_212);
ut213_nn_addition: nn_addition port map( store_weight_426,store_weight_427,sum_213);
ut214_nn_addition: nn_addition port map( store_weight_428,store_weight_429,sum_214);
ut215_nn_addition: nn_addition port map( store_weight_430,store_weight_431,sum_215);
ut216_nn_addition: nn_addition port map( store_weight_432,store_weight_433,sum_216);
ut217_nn_addition: nn_addition port map( store_weight_434,store_weight_435,sum_217);
ut218_nn_addition: nn_addition port map( store_weight_436,store_weight_437,sum_218);
ut219_nn_addition: nn_addition port map( store_weight_438,store_weight_439,sum_219);
ut220_nn_addition: nn_addition port map( store_weight_440,store_weight_441,sum_220);
ut221_nn_addition: nn_addition port map( store_weight_442,store_weight_443,sum_221);
ut222_nn_addition: nn_addition port map( store_weight_444,store_weight_445,sum_222);
ut223_nn_addition: nn_addition port map( store_weight_446,store_weight_447,sum_223);
ut224_nn_addition: nn_addition port map( store_weight_448,store_weight_449,sum_224);
ut225_nn_addition: nn_addition port map( store_weight_450,store_weight_451,sum_225);
ut226_nn_addition: nn_addition port map( store_weight_452,store_weight_453,sum_226);
ut227_nn_addition: nn_addition port map( store_weight_454,store_weight_455,sum_227);
ut228_nn_addition: nn_addition port map( store_weight_456,store_weight_457,sum_228);
ut229_nn_addition: nn_addition port map( store_weight_458,store_weight_459,sum_229);
ut230_nn_addition: nn_addition port map( store_weight_460,store_weight_461,sum_230);
ut231_nn_addition: nn_addition port map( store_weight_462,store_weight_463,sum_231);
ut232_nn_addition: nn_addition port map( store_weight_464,store_weight_465,sum_232);
ut233_nn_addition: nn_addition port map( store_weight_466,store_weight_467,sum_233);
ut234_nn_addition: nn_addition port map( store_weight_468,store_weight_469,sum_234);
ut235_nn_addition: nn_addition port map( store_weight_470,store_weight_471,sum_235);
ut236_nn_addition: nn_addition port map( store_weight_472,store_weight_473,sum_236);
ut237_nn_addition: nn_addition port map( store_weight_474,store_weight_475,sum_237);
ut238_nn_addition: nn_addition port map( store_weight_476,store_weight_477,sum_238);
ut239_nn_addition: nn_addition port map( store_weight_478,store_weight_479,sum_239);
ut240_nn_addition: nn_addition port map( store_weight_480,store_weight_481,sum_240);
ut241_nn_addition: nn_addition port map( store_weight_482,store_weight_483,sum_241);
ut242_nn_addition: nn_addition port map( store_weight_484,store_weight_485,sum_242);
ut243_nn_addition: nn_addition port map( store_weight_486,store_weight_487,sum_243);
ut244_nn_addition: nn_addition port map( store_weight_488,store_weight_489,sum_244);
ut245_nn_addition: nn_addition port map( store_weight_490,store_weight_491,sum_245);
ut246_nn_addition: nn_addition port map( store_weight_492,store_weight_493,sum_246);
ut247_nn_addition: nn_addition port map( store_weight_494,store_weight_495,sum_247);
ut248_nn_addition: nn_addition port map( store_weight_496,store_weight_497,sum_248);
ut249_nn_addition: nn_addition port map( store_weight_498,store_weight_499,sum_249);
ut250_nn_addition: nn_addition port map( store_weight_500,store_weight_501,sum_250);
ut251_nn_addition: nn_addition port map( store_weight_502,store_weight_503,sum_251);
ut252_nn_addition: nn_addition port map( store_weight_504,store_weight_505,sum_252);
ut253_nn_addition: nn_addition port map( store_weight_506,store_weight_507,sum_253);
ut254_nn_addition: nn_addition port map( store_weight_508,store_weight_509,sum_254);
ut255_nn_addition: nn_addition port map( store_weight_510,store_weight_511,sum_255);
ut256_nn_addition: nn_addition port map( store_weight_512,store_weight_513,sum_256);
ut257_nn_addition: nn_addition port map( store_weight_514,store_weight_515,sum_257);
ut258_nn_addition: nn_addition port map( store_weight_516,store_weight_517,sum_258);
ut259_nn_addition: nn_addition port map( store_weight_518,store_weight_519,sum_259);
ut260_nn_addition: nn_addition port map( store_weight_520,store_weight_521,sum_260);
ut261_nn_addition: nn_addition port map( store_weight_522,store_weight_523,sum_261);
ut262_nn_addition: nn_addition port map( store_weight_524,store_weight_525,sum_262);
ut263_nn_addition: nn_addition port map( store_weight_526,store_weight_527,sum_263);
ut264_nn_addition: nn_addition port map( store_weight_528,store_weight_529,sum_264);
ut265_nn_addition: nn_addition port map( store_weight_530,store_weight_531,sum_265);
ut266_nn_addition: nn_addition port map( store_weight_532,store_weight_533,sum_266);
ut267_nn_addition: nn_addition port map( store_weight_534,store_weight_535,sum_267);
ut268_nn_addition: nn_addition port map( store_weight_536,store_weight_537,sum_268);
ut269_nn_addition: nn_addition port map( store_weight_538,store_weight_539,sum_269);
ut270_nn_addition: nn_addition port map( store_weight_540,store_weight_541,sum_270);
ut271_nn_addition: nn_addition port map( store_weight_542,store_weight_543,sum_271);
ut272_nn_addition: nn_addition port map( store_weight_544,store_weight_545,sum_272);
ut273_nn_addition: nn_addition port map( store_weight_546,store_weight_547,sum_273);
ut274_nn_addition: nn_addition port map( store_weight_548,store_weight_549,sum_274);
ut275_nn_addition: nn_addition port map( store_weight_550,store_weight_551,sum_275);
ut276_nn_addition: nn_addition port map( store_weight_552,store_weight_553,sum_276);
ut277_nn_addition: nn_addition port map( store_weight_554,store_weight_555,sum_277);
ut278_nn_addition: nn_addition port map( store_weight_556,store_weight_557,sum_278);
ut279_nn_addition: nn_addition port map( store_weight_558,store_weight_559,sum_279);
ut280_nn_addition: nn_addition port map( store_weight_560,store_weight_561,sum_280);
ut281_nn_addition: nn_addition port map( store_weight_562,store_weight_563,sum_281);
ut282_nn_addition: nn_addition port map( store_weight_564,store_weight_565,sum_282);
ut283_nn_addition: nn_addition port map( store_weight_566,store_weight_567,sum_283);
ut284_nn_addition: nn_addition port map( store_weight_568,store_weight_569,sum_284);
ut285_nn_addition: nn_addition port map( store_weight_570,store_weight_571,sum_285);
ut286_nn_addition: nn_addition port map( store_weight_572,store_weight_573,sum_286);
ut287_nn_addition: nn_addition port map( store_weight_574,store_weight_575,sum_287);
ut288_nn_addition: nn_addition port map( store_weight_576,store_weight_577,sum_288);
ut289_nn_addition: nn_addition port map( store_weight_578,store_weight_579,sum_289);
ut290_nn_addition: nn_addition port map( store_weight_580,store_weight_581,sum_290);
ut291_nn_addition: nn_addition port map( store_weight_582,store_weight_583,sum_291);
ut292_nn_addition: nn_addition port map( store_weight_584,store_weight_585,sum_292);
ut293_nn_addition: nn_addition port map( store_weight_586,store_weight_587,sum_293);
ut294_nn_addition: nn_addition port map( store_weight_588,store_weight_589,sum_294);
ut295_nn_addition: nn_addition port map( store_weight_590,store_weight_591,sum_295);
ut296_nn_addition: nn_addition port map( store_weight_592,store_weight_593,sum_296);
ut297_nn_addition: nn_addition port map( store_weight_594,store_weight_595,sum_297);
ut298_nn_addition: nn_addition port map( store_weight_596,store_weight_597,sum_298);
ut299_nn_addition: nn_addition port map( store_weight_598,store_weight_599,sum_299);
ut300_nn_addition: nn_addition port map( store_weight_600,store_weight_601,sum_300);
ut301_nn_addition: nn_addition port map( store_weight_602,store_weight_603,sum_301);
ut302_nn_addition: nn_addition port map( store_weight_604,store_weight_605,sum_302);
ut303_nn_addition: nn_addition port map( store_weight_606,store_weight_607,sum_303);
ut304_nn_addition: nn_addition port map( store_weight_608,store_weight_609,sum_304);
ut305_nn_addition: nn_addition port map( store_weight_610,store_weight_611,sum_305);
ut306_nn_addition: nn_addition port map( store_weight_612,store_weight_613,sum_306);
ut307_nn_addition: nn_addition port map( store_weight_614,store_weight_615,sum_307);
ut308_nn_addition: nn_addition port map( store_weight_616,store_weight_617,sum_308);
ut309_nn_addition: nn_addition port map( store_weight_618,store_weight_619,sum_309);
ut310_nn_addition: nn_addition port map( store_weight_620,store_weight_621,sum_310);
ut311_nn_addition: nn_addition port map( store_weight_622,store_weight_623,sum_311);
ut312_nn_addition: nn_addition port map( store_weight_624,store_weight_625,sum_312);
ut313_nn_addition: nn_addition port map( store_weight_626,store_weight_627,sum_313);
ut314_nn_addition: nn_addition port map( store_weight_628,store_weight_629,sum_314);
ut315_nn_addition: nn_addition port map( store_weight_630,store_weight_631,sum_315);
ut316_nn_addition: nn_addition port map( store_weight_632,store_weight_633,sum_316);
ut317_nn_addition: nn_addition port map( store_weight_634,store_weight_635,sum_317);
ut318_nn_addition: nn_addition port map( store_weight_636,store_weight_637,sum_318);
ut319_nn_addition: nn_addition port map( store_weight_638,store_weight_639,sum_319);
ut320_nn_addition: nn_addition port map( store_weight_640,store_weight_641,sum_320);
ut321_nn_addition: nn_addition port map( store_weight_642,store_weight_643,sum_321);
ut322_nn_addition: nn_addition port map( store_weight_644,store_weight_645,sum_322);
ut323_nn_addition: nn_addition port map( store_weight_646,store_weight_647,sum_323);
ut324_nn_addition: nn_addition port map( store_weight_648,store_weight_649,sum_324);
ut325_nn_addition: nn_addition port map( store_weight_650,store_weight_651,sum_325);
ut326_nn_addition: nn_addition port map( store_weight_652,store_weight_653,sum_326);
ut327_nn_addition: nn_addition port map( store_weight_654,store_weight_655,sum_327);
ut328_nn_addition: nn_addition port map( store_weight_656,store_weight_657,sum_328);
ut329_nn_addition: nn_addition port map( store_weight_658,store_weight_659,sum_329);
ut330_nn_addition: nn_addition port map( store_weight_660,store_weight_661,sum_330);
ut331_nn_addition: nn_addition port map( store_weight_662,store_weight_663,sum_331);
ut332_nn_addition: nn_addition port map( store_weight_664,store_weight_665,sum_332);
ut333_nn_addition: nn_addition port map( store_weight_666,store_weight_667,sum_333);
ut334_nn_addition: nn_addition port map( store_weight_668,store_weight_669,sum_334);
ut335_nn_addition: nn_addition port map( store_weight_670,store_weight_671,sum_335);
ut336_nn_addition: nn_addition port map( store_weight_672,store_weight_673,sum_336);
ut337_nn_addition: nn_addition port map( store_weight_674,store_weight_675,sum_337);
ut338_nn_addition: nn_addition port map( store_weight_676,store_weight_677,sum_338);
ut339_nn_addition: nn_addition port map( store_weight_678,store_weight_679,sum_339);
ut340_nn_addition: nn_addition port map( store_weight_680,store_weight_681,sum_340);
ut341_nn_addition: nn_addition port map( store_weight_682,store_weight_683,sum_341);
ut342_nn_addition: nn_addition port map( store_weight_684,store_weight_685,sum_342);
ut343_nn_addition: nn_addition port map( store_weight_686,store_weight_687,sum_343);
ut344_nn_addition: nn_addition port map( store_weight_688,store_weight_689,sum_344);
ut345_nn_addition: nn_addition port map( store_weight_690,store_weight_691,sum_345);
ut346_nn_addition: nn_addition port map( store_weight_692,store_weight_693,sum_346);
ut347_nn_addition: nn_addition port map( store_weight_694,store_weight_695,sum_347);
ut348_nn_addition: nn_addition port map( store_weight_696,store_weight_697,sum_348);
ut349_nn_addition: nn_addition port map( store_weight_698,store_weight_699,sum_349);
ut350_nn_addition: nn_addition port map( store_weight_700,store_weight_701,sum_350);
ut351_nn_addition: nn_addition port map( store_weight_702,store_weight_703,sum_351);
ut352_nn_addition: nn_addition port map( store_weight_704,store_weight_705,sum_352);
ut353_nn_addition: nn_addition port map( store_weight_706,store_weight_707,sum_353);
ut354_nn_addition: nn_addition port map( store_weight_708,store_weight_709,sum_354);
ut355_nn_addition: nn_addition port map( store_weight_710,store_weight_711,sum_355);
ut356_nn_addition: nn_addition port map( store_weight_712,store_weight_713,sum_356);
ut357_nn_addition: nn_addition port map( store_weight_714,store_weight_715,sum_357);
ut358_nn_addition: nn_addition port map( store_weight_716,store_weight_717,sum_358);
ut359_nn_addition: nn_addition port map( store_weight_718,store_weight_719,sum_359);
ut360_nn_addition: nn_addition port map( store_weight_720,store_weight_721,sum_360);
ut361_nn_addition: nn_addition port map( store_weight_722,store_weight_723,sum_361);
ut362_nn_addition: nn_addition port map( store_weight_724,store_weight_725,sum_362);
ut363_nn_addition: nn_addition port map( store_weight_726,store_weight_727,sum_363);
ut364_nn_addition: nn_addition port map( store_weight_728,store_weight_729,sum_364);
ut365_nn_addition: nn_addition port map( store_weight_730,store_weight_731,sum_365);
ut366_nn_addition: nn_addition port map( store_weight_732,store_weight_733,sum_366);
ut367_nn_addition: nn_addition port map( store_weight_734,store_weight_735,sum_367);
ut368_nn_addition: nn_addition port map( store_weight_736,store_weight_737,sum_368);
ut369_nn_addition: nn_addition port map( store_weight_738,store_weight_739,sum_369);
ut370_nn_addition: nn_addition port map( store_weight_740,store_weight_741,sum_370);
ut371_nn_addition: nn_addition port map( store_weight_742,store_weight_743,sum_371);
ut372_nn_addition: nn_addition port map( store_weight_744,store_weight_745,sum_372);
ut373_nn_addition: nn_addition port map( store_weight_746,store_weight_747,sum_373);
ut374_nn_addition: nn_addition port map( store_weight_748,store_weight_749,sum_374);
ut375_nn_addition: nn_addition port map( store_weight_750,store_weight_751,sum_375);
ut376_nn_addition: nn_addition port map( store_weight_752,store_weight_753,sum_376);
ut377_nn_addition: nn_addition port map( store_weight_754,store_weight_755,sum_377);
ut378_nn_addition: nn_addition port map( store_weight_756,store_weight_757,sum_378);
ut379_nn_addition: nn_addition port map( store_weight_758,store_weight_759,sum_379);
ut380_nn_addition: nn_addition port map( store_weight_760,store_weight_761,sum_380);
ut381_nn_addition: nn_addition port map( store_weight_762,store_weight_763,sum_381);
ut382_nn_addition: nn_addition port map( store_weight_764,store_weight_765,sum_382);
ut383_nn_addition: nn_addition port map( store_weight_766,store_weight_767,sum_383);
ut384_nn_addition: nn_addition port map( store_weight_768,store_weight_769,sum_384);
ut385_nn_addition: nn_addition port map( store_weight_770,store_weight_771,sum_385);
ut386_nn_addition: nn_addition port map( store_weight_772,store_weight_773,sum_386);
ut387_nn_addition: nn_addition port map( store_weight_774,store_weight_775,sum_387);
ut388_nn_addition: nn_addition port map( store_weight_776,store_weight_777,sum_388);
ut389_nn_addition: nn_addition port map( store_weight_778,store_weight_779,sum_389);
ut390_nn_addition: nn_addition port map( store_weight_780,store_weight_781,sum_390);
ut391_nn_addition: nn_addition port map( store_weight_782,store_weight_783,sum_391);
ut392_nn_addition: nn_addition port map( sum_0,sum_1,sum_392);
ut393_nn_addition: nn_addition port map( sum_2,sum_3,sum_393);
ut394_nn_addition: nn_addition port map( sum_4,sum_5,sum_394);
ut395_nn_addition: nn_addition port map( sum_6,sum_7,sum_395);
ut396_nn_addition: nn_addition port map( sum_8,sum_9,sum_396);
ut397_nn_addition: nn_addition port map( sum_10,sum_11,sum_397);
ut398_nn_addition: nn_addition port map( sum_12,sum_13,sum_398);
ut399_nn_addition: nn_addition port map( sum_14,sum_15,sum_399);
ut400_nn_addition: nn_addition port map( sum_16,sum_17,sum_400);
ut401_nn_addition: nn_addition port map( sum_18,sum_19,sum_401);
ut402_nn_addition: nn_addition port map( sum_20,sum_21,sum_402);
ut403_nn_addition: nn_addition port map( sum_22,sum_23,sum_403);
ut404_nn_addition: nn_addition port map( sum_24,sum_25,sum_404);
ut405_nn_addition: nn_addition port map( sum_26,sum_27,sum_405);
ut406_nn_addition: nn_addition port map( sum_28,sum_29,sum_406);
ut407_nn_addition: nn_addition port map( sum_30,sum_31,sum_407);
ut408_nn_addition: nn_addition port map( sum_32,sum_33,sum_408);
ut409_nn_addition: nn_addition port map( sum_34,sum_35,sum_409);
ut410_nn_addition: nn_addition port map( sum_36,sum_37,sum_410);
ut411_nn_addition: nn_addition port map( sum_38,sum_39,sum_411);
ut412_nn_addition: nn_addition port map( sum_40,sum_41,sum_412);
ut413_nn_addition: nn_addition port map( sum_42,sum_43,sum_413);
ut414_nn_addition: nn_addition port map( sum_44,sum_45,sum_414);
ut415_nn_addition: nn_addition port map( sum_46,sum_47,sum_415);
ut416_nn_addition: nn_addition port map( sum_48,sum_49,sum_416);
ut417_nn_addition: nn_addition port map( sum_50,sum_51,sum_417);
ut418_nn_addition: nn_addition port map( sum_52,sum_53,sum_418);
ut419_nn_addition: nn_addition port map( sum_54,sum_55,sum_419);
ut420_nn_addition: nn_addition port map( sum_56,sum_57,sum_420);
ut421_nn_addition: nn_addition port map( sum_58,sum_59,sum_421);
ut422_nn_addition: nn_addition port map( sum_60,sum_61,sum_422);
ut423_nn_addition: nn_addition port map( sum_62,sum_63,sum_423);
ut424_nn_addition: nn_addition port map( sum_64,sum_65,sum_424);
ut425_nn_addition: nn_addition port map( sum_66,sum_67,sum_425);
ut426_nn_addition: nn_addition port map( sum_68,sum_69,sum_426);
ut427_nn_addition: nn_addition port map( sum_70,sum_71,sum_427);
ut428_nn_addition: nn_addition port map( sum_72,sum_73,sum_428);
ut429_nn_addition: nn_addition port map( sum_74,sum_75,sum_429);
ut430_nn_addition: nn_addition port map( sum_76,sum_77,sum_430);
ut431_nn_addition: nn_addition port map( sum_78,sum_79,sum_431);
ut432_nn_addition: nn_addition port map( sum_80,sum_81,sum_432);
ut433_nn_addition: nn_addition port map( sum_82,sum_83,sum_433);
ut434_nn_addition: nn_addition port map( sum_84,sum_85,sum_434);
ut435_nn_addition: nn_addition port map( sum_86,sum_87,sum_435);
ut436_nn_addition: nn_addition port map( sum_88,sum_89,sum_436);
ut437_nn_addition: nn_addition port map( sum_90,sum_91,sum_437);
ut438_nn_addition: nn_addition port map( sum_92,sum_93,sum_438);
ut439_nn_addition: nn_addition port map( sum_94,sum_95,sum_439);
ut440_nn_addition: nn_addition port map( sum_96,sum_97,sum_440);
ut441_nn_addition: nn_addition port map( sum_98,sum_99,sum_441);
ut442_nn_addition: nn_addition port map( sum_100,sum_101,sum_442);
ut443_nn_addition: nn_addition port map( sum_102,sum_103,sum_443);
ut444_nn_addition: nn_addition port map( sum_104,sum_105,sum_444);
ut445_nn_addition: nn_addition port map( sum_106,sum_107,sum_445);
ut446_nn_addition: nn_addition port map( sum_108,sum_109,sum_446);
ut447_nn_addition: nn_addition port map( sum_110,sum_111,sum_447);
ut448_nn_addition: nn_addition port map( sum_112,sum_113,sum_448);
ut449_nn_addition: nn_addition port map( sum_114,sum_115,sum_449);
ut450_nn_addition: nn_addition port map( sum_116,sum_117,sum_450);
ut451_nn_addition: nn_addition port map( sum_118,sum_119,sum_451);
ut452_nn_addition: nn_addition port map( sum_120,sum_121,sum_452);
ut453_nn_addition: nn_addition port map( sum_122,sum_123,sum_453);
ut454_nn_addition: nn_addition port map( sum_124,sum_125,sum_454);
ut455_nn_addition: nn_addition port map( sum_126,sum_127,sum_455);
ut456_nn_addition: nn_addition port map( sum_128,sum_129,sum_456);
ut457_nn_addition: nn_addition port map( sum_130,sum_131,sum_457);
ut458_nn_addition: nn_addition port map( sum_132,sum_133,sum_458);
ut459_nn_addition: nn_addition port map( sum_134,sum_135,sum_459);
ut460_nn_addition: nn_addition port map( sum_136,sum_137,sum_460);
ut461_nn_addition: nn_addition port map( sum_138,sum_139,sum_461);
ut462_nn_addition: nn_addition port map( sum_140,sum_141,sum_462);
ut463_nn_addition: nn_addition port map( sum_142,sum_143,sum_463);
ut464_nn_addition: nn_addition port map( sum_144,sum_145,sum_464);
ut465_nn_addition: nn_addition port map( sum_146,sum_147,sum_465);
ut466_nn_addition: nn_addition port map( sum_148,sum_149,sum_466);
ut467_nn_addition: nn_addition port map( sum_150,sum_151,sum_467);
ut468_nn_addition: nn_addition port map( sum_152,sum_153,sum_468);
ut469_nn_addition: nn_addition port map( sum_154,sum_155,sum_469);
ut470_nn_addition: nn_addition port map( sum_156,sum_157,sum_470);
ut471_nn_addition: nn_addition port map( sum_158,sum_159,sum_471);
ut472_nn_addition: nn_addition port map( sum_160,sum_161,sum_472);
ut473_nn_addition: nn_addition port map( sum_162,sum_163,sum_473);
ut474_nn_addition: nn_addition port map( sum_164,sum_165,sum_474);
ut475_nn_addition: nn_addition port map( sum_166,sum_167,sum_475);
ut476_nn_addition: nn_addition port map( sum_168,sum_169,sum_476);
ut477_nn_addition: nn_addition port map( sum_170,sum_171,sum_477);
ut478_nn_addition: nn_addition port map( sum_172,sum_173,sum_478);
ut479_nn_addition: nn_addition port map( sum_174,sum_175,sum_479);
ut480_nn_addition: nn_addition port map( sum_176,sum_177,sum_480);
ut481_nn_addition: nn_addition port map( sum_178,sum_179,sum_481);
ut482_nn_addition: nn_addition port map( sum_180,sum_181,sum_482);
ut483_nn_addition: nn_addition port map( sum_182,sum_183,sum_483);
ut484_nn_addition: nn_addition port map( sum_184,sum_185,sum_484);
ut485_nn_addition: nn_addition port map( sum_186,sum_187,sum_485);
ut486_nn_addition: nn_addition port map( sum_188,sum_189,sum_486);
ut487_nn_addition: nn_addition port map( sum_190,sum_191,sum_487);
ut488_nn_addition: nn_addition port map( sum_192,sum_193,sum_488);
ut489_nn_addition: nn_addition port map( sum_194,sum_195,sum_489);
ut490_nn_addition: nn_addition port map( sum_196,sum_197,sum_490);
ut491_nn_addition: nn_addition port map( sum_198,sum_199,sum_491);
ut492_nn_addition: nn_addition port map( sum_200,sum_201,sum_492);
ut493_nn_addition: nn_addition port map( sum_202,sum_203,sum_493);
ut494_nn_addition: nn_addition port map( sum_204,sum_205,sum_494);
ut495_nn_addition: nn_addition port map( sum_206,sum_207,sum_495);
ut496_nn_addition: nn_addition port map( sum_208,sum_209,sum_496);
ut497_nn_addition: nn_addition port map( sum_210,sum_211,sum_497);
ut498_nn_addition: nn_addition port map( sum_212,sum_213,sum_498);
ut499_nn_addition: nn_addition port map( sum_214,sum_215,sum_499);
ut500_nn_addition: nn_addition port map( sum_216,sum_217,sum_500);
ut501_nn_addition: nn_addition port map( sum_218,sum_219,sum_501);
ut502_nn_addition: nn_addition port map( sum_220,sum_221,sum_502);
ut503_nn_addition: nn_addition port map( sum_222,sum_223,sum_503);
ut504_nn_addition: nn_addition port map( sum_224,sum_225,sum_504);
ut505_nn_addition: nn_addition port map( sum_226,sum_227,sum_505);
ut506_nn_addition: nn_addition port map( sum_228,sum_229,sum_506);
ut507_nn_addition: nn_addition port map( sum_230,sum_231,sum_507);
ut508_nn_addition: nn_addition port map( sum_232,sum_233,sum_508);
ut509_nn_addition: nn_addition port map( sum_234,sum_235,sum_509);
ut510_nn_addition: nn_addition port map( sum_236,sum_237,sum_510);
ut511_nn_addition: nn_addition port map( sum_238,sum_239,sum_511);
ut512_nn_addition: nn_addition port map( sum_240,sum_241,sum_512);
ut513_nn_addition: nn_addition port map( sum_242,sum_243,sum_513);
ut514_nn_addition: nn_addition port map( sum_244,sum_245,sum_514);
ut515_nn_addition: nn_addition port map( sum_246,sum_247,sum_515);
ut516_nn_addition: nn_addition port map( sum_248,sum_249,sum_516);
ut517_nn_addition: nn_addition port map( sum_250,sum_251,sum_517);
ut518_nn_addition: nn_addition port map( sum_252,sum_253,sum_518);
ut519_nn_addition: nn_addition port map( sum_254,sum_255,sum_519);
ut520_nn_addition: nn_addition port map( sum_256,sum_257,sum_520);
ut521_nn_addition: nn_addition port map( sum_258,sum_259,sum_521);
ut522_nn_addition: nn_addition port map( sum_260,sum_261,sum_522);
ut523_nn_addition: nn_addition port map( sum_262,sum_263,sum_523);
ut524_nn_addition: nn_addition port map( sum_264,sum_265,sum_524);
ut525_nn_addition: nn_addition port map( sum_266,sum_267,sum_525);
ut526_nn_addition: nn_addition port map( sum_268,sum_269,sum_526);
ut527_nn_addition: nn_addition port map( sum_270,sum_271,sum_527);
ut528_nn_addition: nn_addition port map( sum_272,sum_273,sum_528);
ut529_nn_addition: nn_addition port map( sum_274,sum_275,sum_529);
ut530_nn_addition: nn_addition port map( sum_276,sum_277,sum_530);
ut531_nn_addition: nn_addition port map( sum_278,sum_279,sum_531);
ut532_nn_addition: nn_addition port map( sum_280,sum_281,sum_532);
ut533_nn_addition: nn_addition port map( sum_282,sum_283,sum_533);
ut534_nn_addition: nn_addition port map( sum_284,sum_285,sum_534);
ut535_nn_addition: nn_addition port map( sum_286,sum_287,sum_535);
ut536_nn_addition: nn_addition port map( sum_288,sum_289,sum_536);
ut537_nn_addition: nn_addition port map( sum_290,sum_291,sum_537);
ut538_nn_addition: nn_addition port map( sum_292,sum_293,sum_538);
ut539_nn_addition: nn_addition port map( sum_294,sum_295,sum_539);
ut540_nn_addition: nn_addition port map( sum_296,sum_297,sum_540);
ut541_nn_addition: nn_addition port map( sum_298,sum_299,sum_541);
ut542_nn_addition: nn_addition port map( sum_300,sum_301,sum_542);
ut543_nn_addition: nn_addition port map( sum_302,sum_303,sum_543);
ut544_nn_addition: nn_addition port map( sum_304,sum_305,sum_544);
ut545_nn_addition: nn_addition port map( sum_306,sum_307,sum_545);
ut546_nn_addition: nn_addition port map( sum_308,sum_309,sum_546);
ut547_nn_addition: nn_addition port map( sum_310,sum_311,sum_547);
ut548_nn_addition: nn_addition port map( sum_312,sum_313,sum_548);
ut549_nn_addition: nn_addition port map( sum_314,sum_315,sum_549);
ut550_nn_addition: nn_addition port map( sum_316,sum_317,sum_550);
ut551_nn_addition: nn_addition port map( sum_318,sum_319,sum_551);
ut552_nn_addition: nn_addition port map( sum_320,sum_321,sum_552);
ut553_nn_addition: nn_addition port map( sum_322,sum_323,sum_553);
ut554_nn_addition: nn_addition port map( sum_324,sum_325,sum_554);
ut555_nn_addition: nn_addition port map( sum_326,sum_327,sum_555);
ut556_nn_addition: nn_addition port map( sum_328,sum_329,sum_556);
ut557_nn_addition: nn_addition port map( sum_330,sum_331,sum_557);
ut558_nn_addition: nn_addition port map( sum_332,sum_333,sum_558);
ut559_nn_addition: nn_addition port map( sum_334,sum_335,sum_559);
ut560_nn_addition: nn_addition port map( sum_336,sum_337,sum_560);
ut561_nn_addition: nn_addition port map( sum_338,sum_339,sum_561);
ut562_nn_addition: nn_addition port map( sum_340,sum_341,sum_562);
ut563_nn_addition: nn_addition port map( sum_342,sum_343,sum_563);
ut564_nn_addition: nn_addition port map( sum_344,sum_345,sum_564);
ut565_nn_addition: nn_addition port map( sum_346,sum_347,sum_565);
ut566_nn_addition: nn_addition port map( sum_348,sum_349,sum_566);
ut567_nn_addition: nn_addition port map( sum_350,sum_351,sum_567);
ut568_nn_addition: nn_addition port map( sum_352,sum_353,sum_568);
ut569_nn_addition: nn_addition port map( sum_354,sum_355,sum_569);
ut570_nn_addition: nn_addition port map( sum_356,sum_357,sum_570);
ut571_nn_addition: nn_addition port map( sum_358,sum_359,sum_571);
ut572_nn_addition: nn_addition port map( sum_360,sum_361,sum_572);
ut573_nn_addition: nn_addition port map( sum_362,sum_363,sum_573);
ut574_nn_addition: nn_addition port map( sum_364,sum_365,sum_574);
ut575_nn_addition: nn_addition port map( sum_366,sum_367,sum_575);
ut576_nn_addition: nn_addition port map( sum_368,sum_369,sum_576);
ut577_nn_addition: nn_addition port map( sum_370,sum_371,sum_577);
ut578_nn_addition: nn_addition port map( sum_372,sum_373,sum_578);
ut579_nn_addition: nn_addition port map( sum_374,sum_375,sum_579);
ut580_nn_addition: nn_addition port map( sum_376,sum_377,sum_580);
ut581_nn_addition: nn_addition port map( sum_378,sum_379,sum_581);
ut582_nn_addition: nn_addition port map( sum_380,sum_381,sum_582);
ut583_nn_addition: nn_addition port map( sum_382,sum_383,sum_583);
ut584_nn_addition: nn_addition port map( sum_384,sum_385,sum_584);
ut585_nn_addition: nn_addition port map( sum_386,sum_387,sum_585);
ut586_nn_addition: nn_addition port map( sum_388,sum_389,sum_586);
ut587_nn_addition: nn_addition port map( sum_390,sum_391,sum_587);
ut588_nn_addition: nn_addition port map( sum_392,sum_393,sum_588);
ut589_nn_addition: nn_addition port map( sum_394,sum_395,sum_589);
ut590_nn_addition: nn_addition port map( sum_396,sum_397,sum_590);
ut591_nn_addition: nn_addition port map( sum_398,sum_399,sum_591);
ut592_nn_addition: nn_addition port map( sum_400,sum_401,sum_592);
ut593_nn_addition: nn_addition port map( sum_402,sum_403,sum_593);
ut594_nn_addition: nn_addition port map( sum_404,sum_405,sum_594);
ut595_nn_addition: nn_addition port map( sum_406,sum_407,sum_595);
ut596_nn_addition: nn_addition port map( sum_408,sum_409,sum_596);
ut597_nn_addition: nn_addition port map( sum_410,sum_411,sum_597);
ut598_nn_addition: nn_addition port map( sum_412,sum_413,sum_598);
ut599_nn_addition: nn_addition port map( sum_414,sum_415,sum_599);
ut600_nn_addition: nn_addition port map( sum_416,sum_417,sum_600);
ut601_nn_addition: nn_addition port map( sum_418,sum_419,sum_601);
ut602_nn_addition: nn_addition port map( sum_420,sum_421,sum_602);
ut603_nn_addition: nn_addition port map( sum_422,sum_423,sum_603);
ut604_nn_addition: nn_addition port map( sum_424,sum_425,sum_604);
ut605_nn_addition: nn_addition port map( sum_426,sum_427,sum_605);
ut606_nn_addition: nn_addition port map( sum_428,sum_429,sum_606);
ut607_nn_addition: nn_addition port map( sum_430,sum_431,sum_607);
ut608_nn_addition: nn_addition port map( sum_432,sum_433,sum_608);
ut609_nn_addition: nn_addition port map( sum_434,sum_435,sum_609);
ut610_nn_addition: nn_addition port map( sum_436,sum_437,sum_610);
ut611_nn_addition: nn_addition port map( sum_438,sum_439,sum_611);
ut612_nn_addition: nn_addition port map( sum_440,sum_441,sum_612);
ut613_nn_addition: nn_addition port map( sum_442,sum_443,sum_613);
ut614_nn_addition: nn_addition port map( sum_444,sum_445,sum_614);
ut615_nn_addition: nn_addition port map( sum_446,sum_447,sum_615);
ut616_nn_addition: nn_addition port map( sum_448,sum_449,sum_616);
ut617_nn_addition: nn_addition port map( sum_450,sum_451,sum_617);
ut618_nn_addition: nn_addition port map( sum_452,sum_453,sum_618);
ut619_nn_addition: nn_addition port map( sum_454,sum_455,sum_619);
ut620_nn_addition: nn_addition port map( sum_456,sum_457,sum_620);
ut621_nn_addition: nn_addition port map( sum_458,sum_459,sum_621);
ut622_nn_addition: nn_addition port map( sum_460,sum_461,sum_622);
ut623_nn_addition: nn_addition port map( sum_462,sum_463,sum_623);
ut624_nn_addition: nn_addition port map( sum_464,sum_465,sum_624);
ut625_nn_addition: nn_addition port map( sum_466,sum_467,sum_625);
ut626_nn_addition: nn_addition port map( sum_468,sum_469,sum_626);
ut627_nn_addition: nn_addition port map( sum_470,sum_471,sum_627);
ut628_nn_addition: nn_addition port map( sum_472,sum_473,sum_628);
ut629_nn_addition: nn_addition port map( sum_474,sum_475,sum_629);
ut630_nn_addition: nn_addition port map( sum_476,sum_477,sum_630);
ut631_nn_addition: nn_addition port map( sum_478,sum_479,sum_631);
ut632_nn_addition: nn_addition port map( sum_480,sum_481,sum_632);
ut633_nn_addition: nn_addition port map( sum_482,sum_483,sum_633);
ut634_nn_addition: nn_addition port map( sum_484,sum_485,sum_634);
ut635_nn_addition: nn_addition port map( sum_486,sum_487,sum_635);
ut636_nn_addition: nn_addition port map( sum_488,sum_489,sum_636);
ut637_nn_addition: nn_addition port map( sum_490,sum_491,sum_637);
ut638_nn_addition: nn_addition port map( sum_492,sum_493,sum_638);
ut639_nn_addition: nn_addition port map( sum_494,sum_495,sum_639);
ut640_nn_addition: nn_addition port map( sum_496,sum_497,sum_640);
ut641_nn_addition: nn_addition port map( sum_498,sum_499,sum_641);
ut642_nn_addition: nn_addition port map( sum_500,sum_501,sum_642);
ut643_nn_addition: nn_addition port map( sum_502,sum_503,sum_643);
ut644_nn_addition: nn_addition port map( sum_504,sum_505,sum_644);
ut645_nn_addition: nn_addition port map( sum_506,sum_507,sum_645);
ut646_nn_addition: nn_addition port map( sum_508,sum_509,sum_646);
ut647_nn_addition: nn_addition port map( sum_510,sum_511,sum_647);
ut648_nn_addition: nn_addition port map( sum_512,sum_513,sum_648);
ut649_nn_addition: nn_addition port map( sum_514,sum_515,sum_649);
ut650_nn_addition: nn_addition port map( sum_516,sum_517,sum_650);
ut651_nn_addition: nn_addition port map( sum_518,sum_519,sum_651);
ut652_nn_addition: nn_addition port map( sum_520,sum_521,sum_652);
ut653_nn_addition: nn_addition port map( sum_522,sum_523,sum_653);
ut654_nn_addition: nn_addition port map( sum_524,sum_525,sum_654);
ut655_nn_addition: nn_addition port map( sum_526,sum_527,sum_655);
ut656_nn_addition: nn_addition port map( sum_528,sum_529,sum_656);
ut657_nn_addition: nn_addition port map( sum_530,sum_531,sum_657);
ut658_nn_addition: nn_addition port map( sum_532,sum_533,sum_658);
ut659_nn_addition: nn_addition port map( sum_534,sum_535,sum_659);
ut660_nn_addition: nn_addition port map( sum_536,sum_537,sum_660);
ut661_nn_addition: nn_addition port map( sum_538,sum_539,sum_661);
ut662_nn_addition: nn_addition port map( sum_540,sum_541,sum_662);
ut663_nn_addition: nn_addition port map( sum_542,sum_543,sum_663);
ut664_nn_addition: nn_addition port map( sum_544,sum_545,sum_664);
ut665_nn_addition: nn_addition port map( sum_546,sum_547,sum_665);
ut666_nn_addition: nn_addition port map( sum_548,sum_549,sum_666);
ut667_nn_addition: nn_addition port map( sum_550,sum_551,sum_667);
ut668_nn_addition: nn_addition port map( sum_552,sum_553,sum_668);
ut669_nn_addition: nn_addition port map( sum_554,sum_555,sum_669);
ut670_nn_addition: nn_addition port map( sum_556,sum_557,sum_670);
ut671_nn_addition: nn_addition port map( sum_558,sum_559,sum_671);
ut672_nn_addition: nn_addition port map( sum_560,sum_561,sum_672);
ut673_nn_addition: nn_addition port map( sum_562,sum_563,sum_673);
ut674_nn_addition: nn_addition port map( sum_564,sum_565,sum_674);
ut675_nn_addition: nn_addition port map( sum_566,sum_567,sum_675);
ut676_nn_addition: nn_addition port map( sum_568,sum_569,sum_676);
ut677_nn_addition: nn_addition port map( sum_570,sum_571,sum_677);
ut678_nn_addition: nn_addition port map( sum_572,sum_573,sum_678);
ut679_nn_addition: nn_addition port map( sum_574,sum_575,sum_679);
ut680_nn_addition: nn_addition port map( sum_576,sum_577,sum_680);
ut681_nn_addition: nn_addition port map( sum_578,sum_579,sum_681);
ut682_nn_addition: nn_addition port map( sum_580,sum_581,sum_682);
ut683_nn_addition: nn_addition port map( sum_582,sum_583,sum_683);
ut684_nn_addition: nn_addition port map( sum_584,sum_585,sum_684);
ut685_nn_addition: nn_addition port map( sum_586,sum_587,sum_685);
ut686_nn_addition: nn_addition port map( sum_588,sum_589,sum_686);
ut687_nn_addition: nn_addition port map( sum_590,sum_591,sum_687);
ut688_nn_addition: nn_addition port map( sum_592,sum_593,sum_688);
ut689_nn_addition: nn_addition port map( sum_594,sum_595,sum_689);
ut690_nn_addition: nn_addition port map( sum_596,sum_597,sum_690);
ut691_nn_addition: nn_addition port map( sum_598,sum_599,sum_691);
ut692_nn_addition: nn_addition port map( sum_600,sum_601,sum_692);
ut693_nn_addition: nn_addition port map( sum_602,sum_603,sum_693);
ut694_nn_addition: nn_addition port map( sum_604,sum_605,sum_694);
ut695_nn_addition: nn_addition port map( sum_606,sum_607,sum_695);
ut696_nn_addition: nn_addition port map( sum_608,sum_609,sum_696);
ut697_nn_addition: nn_addition port map( sum_610,sum_611,sum_697);
ut698_nn_addition: nn_addition port map( sum_612,sum_613,sum_698);
ut699_nn_addition: nn_addition port map( sum_614,sum_615,sum_699);
ut700_nn_addition: nn_addition port map( sum_616,sum_617,sum_700);
ut701_nn_addition: nn_addition port map( sum_618,sum_619,sum_701);
ut702_nn_addition: nn_addition port map( sum_620,sum_621,sum_702);
ut703_nn_addition: nn_addition port map( sum_622,sum_623,sum_703);
ut704_nn_addition: nn_addition port map( sum_624,sum_625,sum_704);
ut705_nn_addition: nn_addition port map( sum_626,sum_627,sum_705);
ut706_nn_addition: nn_addition port map( sum_628,sum_629,sum_706);
ut707_nn_addition: nn_addition port map( sum_630,sum_631,sum_707);
ut708_nn_addition: nn_addition port map( sum_632,sum_633,sum_708);
ut709_nn_addition: nn_addition port map( sum_634,sum_635,sum_709);
ut710_nn_addition: nn_addition port map( sum_636,sum_637,sum_710);
ut711_nn_addition: nn_addition port map( sum_638,sum_639,sum_711);
ut712_nn_addition: nn_addition port map( sum_640,sum_641,sum_712);
ut713_nn_addition: nn_addition port map( sum_642,sum_643,sum_713);
ut714_nn_addition: nn_addition port map( sum_644,sum_645,sum_714);
ut715_nn_addition: nn_addition port map( sum_646,sum_647,sum_715);
ut716_nn_addition: nn_addition port map( sum_648,sum_649,sum_716);
ut717_nn_addition: nn_addition port map( sum_650,sum_651,sum_717);
ut718_nn_addition: nn_addition port map( sum_652,sum_653,sum_718);
ut719_nn_addition: nn_addition port map( sum_654,sum_655,sum_719);
ut720_nn_addition: nn_addition port map( sum_656,sum_657,sum_720);
ut721_nn_addition: nn_addition port map( sum_658,sum_659,sum_721);
ut722_nn_addition: nn_addition port map( sum_660,sum_661,sum_722);
ut723_nn_addition: nn_addition port map( sum_662,sum_663,sum_723);
ut724_nn_addition: nn_addition port map( sum_664,sum_665,sum_724);
ut725_nn_addition: nn_addition port map( sum_666,sum_667,sum_725);
ut726_nn_addition: nn_addition port map( sum_668,sum_669,sum_726);
ut727_nn_addition: nn_addition port map( sum_670,sum_671,sum_727);
ut728_nn_addition: nn_addition port map( sum_672,sum_673,sum_728);
ut729_nn_addition: nn_addition port map( sum_674,sum_675,sum_729);
ut730_nn_addition: nn_addition port map( sum_676,sum_677,sum_730);
ut731_nn_addition: nn_addition port map( sum_678,sum_679,sum_731);
ut732_nn_addition: nn_addition port map( sum_680,sum_681,sum_732);
ut733_nn_addition: nn_addition port map( sum_682,sum_683,sum_733);
ut734_nn_addition: nn_addition port map( sum_684,sum_685,sum_734);
ut735_nn_addition: nn_addition port map( sum_686,sum_687,sum_735);
ut736_nn_addition: nn_addition port map( sum_688,sum_689,sum_736);
ut737_nn_addition: nn_addition port map( sum_690,sum_691,sum_737);
ut738_nn_addition: nn_addition port map( sum_692,sum_693,sum_738);
ut739_nn_addition: nn_addition port map( sum_694,sum_695,sum_739);
ut740_nn_addition: nn_addition port map( sum_696,sum_697,sum_740);
ut741_nn_addition: nn_addition port map( sum_698,sum_699,sum_741);
ut742_nn_addition: nn_addition port map( sum_700,sum_701,sum_742);
ut743_nn_addition: nn_addition port map( sum_702,sum_703,sum_743);
ut744_nn_addition: nn_addition port map( sum_704,sum_705,sum_744);
ut745_nn_addition: nn_addition port map( sum_706,sum_707,sum_745);
ut746_nn_addition: nn_addition port map( sum_708,sum_709,sum_746);
ut747_nn_addition: nn_addition port map( sum_710,sum_711,sum_747);
ut748_nn_addition: nn_addition port map( sum_712,sum_713,sum_748);
ut749_nn_addition: nn_addition port map( sum_714,sum_715,sum_749);
ut750_nn_addition: nn_addition port map( sum_716,sum_717,sum_750);
ut751_nn_addition: nn_addition port map( sum_718,sum_719,sum_751);
ut752_nn_addition: nn_addition port map( sum_720,sum_721,sum_752);
ut753_nn_addition: nn_addition port map( sum_722,sum_723,sum_753);
ut754_nn_addition: nn_addition port map( sum_724,sum_725,sum_754);
ut755_nn_addition: nn_addition port map( sum_726,sum_727,sum_755);
ut756_nn_addition: nn_addition port map( sum_728,sum_729,sum_756);
ut757_nn_addition: nn_addition port map( sum_730,sum_731,sum_757);
ut758_nn_addition: nn_addition port map( sum_732,sum_733,sum_758);
ut759_nn_addition: nn_addition port map( sum_734,sum_735,sum_759);
ut760_nn_addition: nn_addition port map( sum_736,sum_737,sum_760);
ut761_nn_addition: nn_addition port map( sum_738,sum_739,sum_761);
ut762_nn_addition: nn_addition port map( sum_740,sum_741,sum_762);
ut763_nn_addition: nn_addition port map( sum_742,sum_743,sum_763);
ut764_nn_addition: nn_addition port map( sum_744,sum_745,sum_764);
ut765_nn_addition: nn_addition port map( sum_746,sum_747,sum_765);
ut766_nn_addition: nn_addition port map( sum_748,sum_749,sum_766);
ut767_nn_addition: nn_addition port map( sum_750,sum_751,sum_767);
ut768_nn_addition: nn_addition port map( sum_752,sum_753,sum_768);
ut769_nn_addition: nn_addition port map( sum_754,sum_755,sum_769);
ut770_nn_addition: nn_addition port map( sum_756,sum_757,sum_770);
ut771_nn_addition: nn_addition port map( sum_758,sum_759,sum_771);
ut772_nn_addition: nn_addition port map( sum_760,sum_761,sum_772);
ut773_nn_addition: nn_addition port map( sum_762,sum_763,sum_773);
ut774_nn_addition: nn_addition port map( sum_764,sum_765,sum_774);
ut775_nn_addition: nn_addition port map( sum_766,sum_767,sum_775);
ut776_nn_addition: nn_addition port map( sum_768,sum_769,sum_776);
ut777_nn_addition: nn_addition port map( sum_770,sum_771,sum_777);
ut778_nn_addition: nn_addition port map( sum_772,sum_773,sum_778);
ut779_nn_addition: nn_addition port map( sum_774,sum_775,sum_779);
ut780_nn_addition: nn_addition port map( sum_776,sum_777,sum_780);
ut781_nn_addition: nn_addition port map( sum_778,sum_779,sum_781);
ut782_nn_addition: nn_addition port map( sum_780,sum_781,sum_782);
ut784_nn_addition: nn_addition port map( biases,sum_782 ,store_value);
ut1_sigmoid: sigmoid port map( to_integer(unsigned(store_value)),y_3);
end Behavioral;