library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_2 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_2;

architecture syn of ram_2 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"0000000000000111","1000000000001111","0000000000010000","1000000000000101","0000000000010101","1000000000001010","1000000000000011","0000000000001001","0000000000000011","1000000000010001","1000000000001100","1000000000000100","0000000001000011","0000000001000100","1000000000110011","1000000000001000","1000000000010100","1000000000010101","1000000000001100","1000000000001000","1000000000000100","1000000000000101","0000000000010000","0000000000001000","1000000000000110","1000000000000010","1000000000010011","1000000000000011","0000000000010010","1000000000010001","1000000000000000","0000000000000001","0000000000101011","0000000000010101","0000000010100111","0000000010001000","0000000000100010","0000000000111011","0000000011001011","0000000001111000","0000000001111100","0000000010001110","0000000100001101","0000000100010001","0000000010111001","0000000000001000","0000000011010011","0000000100010001","0000000011010000","0000000011000100","0000000010110101","0000000000101011","1000000000010010","1000000000000100","0000000000001001","0000000000001100","1000000000001001","1000000000001000","0000000000010000","1000000000100101","1000000000101000","1000000000101101","1000000001011100","0000000001101110","0000000000110010","0000000010011000","0000000010011010","0000000010100100","0000000100011001","0000000100110110","0000000100101101","0000000100101101","0000000100100110","0000000000111100","0000000000011000","1000000000010010","1000000000001111","0000000011111100","0000000001000001","0000000000010001","0000000000011111","1000000001101000","1000000000010011","1000000000010100","1000000000000100","1000000000010100","0000000010000010","1000000000111000","1000000010100111","0000000000010010","0000000010001001","1000000000100000","1000000100111101","1000000000110011","1000000001011010","1000000011000101","1000000001001010","1000000000110001","1000000010011111","1000000001011010","1000000001000010","1000000010001001","1000000000100000","0000000000111001","1000000000001111","1000000000100101","0000000011000001","0000000000111000","1000000001101000","1000000000101000","1000000001011011","0000000000000011","0000000000000110","1000000000000011","0000000001001011","1000000010100010","0000000000101110","1000000001110111","1000000001100000","1000000001000101","1000000000110111","1000000001001111","1000000000101101","1000000100001100","1000000011100011","1000000011100000","1000000010101001","1000000001111001","1000000000001100","0000000000100110","0000000000001001","0000000000011101","0000000001100110","1000000000010001","0000000001101110","0000000011001111","1000000000000101","1000000000001010","1000000011011000","0000000000100111","0000000000000101","0000000000000100","0000000100111000","1000000010011100","0000000000100010","1000000001000001","0000000000111001","0000000001011001","0000000000011101","1000000001010101","1000000011000101","1000000010111010","1000000010011001","1000000100010110","1000000010110110","1000000001100100","1000000010001111","1000000010001001","1000000001001000","1000000000000111","0000000000000110","0000000000100000","0000000001100001","0000000000100001","0000000010011101","1000000000100110","1000000001101100","0000000001101100","1000000000001001","1000000000011010","1000000010011011","1000000001010010","0000000000001010","1000000100001110","1000000010100011","1000000010011111","1000000011101011","1000000010010100","1000000010001111","1000000010010110","1000000010001011","1000000001111110","1000000000011100","1000000000100110","1000000001011110","1000000001000001","1000000000111111","1000000000101111","1000000001000101","0000000000001000","0000000000101101","0000000000100100","0000000010100010","0000000001010010","1000000010000110","0000000001100110","0000000000111000","1000000001111110","1000000001100011","0000000000000111","1000000001100100","1000000010101100","1000000011011111","1000000010001110","1000000011100101","1000000001000010","1000000001101000","1000000000111110","1000000001100111","1000000000101001","0000000000011001","1000000000100110","1000000000100011","1000000000101111","1000000001111010","1000000000010101","0000000001000000","0000000000000110","0000000000101000","0000000000110011","0000000000110010","1000000100100010","0000000000001101","0000000000011110","1000000001110111","1000000001111100","1000000001001110","0000000000100011","0000000000010100","1000000001111010","1000000000101110","1000000001000111","1000000001100100","1000000000110101","1000000001000000","1000000011010011","1000000001110110","1000000001101000","1000000001001001","1000000001010011","1000000100000010","1000000010100001","1000000001110100","1000000010010010","1000000001101010","1000000001010011","1000000001001010","1000000001011111","1000000010011101","1000000011100100","1000000000011110","1000000010110110","0000000001001011","0000000101101101","0000000000011010","1000000000001110","1000000001010100","1000000100000000","1000000010101011","1000000001100010","1000000010101001","1000000010101010","1000000001110101","1000000001110000","1000000001000011","1000000001000000","0000000000100100","0000000000101101","1000000010001000","1000000101001111","1000000011100001","1000000010111101","1000000011001000","1000000001001001","1000000001110101","1000000011100100","1000000011110110","1000000100000000","1000000001111110","0000000001000110","0000000000111011","0000000111110010","0000000001000001","0000000000001010","1000000010001011","1000000011000100","1000000010111000","1000000000110010","0000000000010101","1000000000100111","1000000000001101","0000000000011100","0000000000110011","0000000001000000","0000000010100000","0000000010111111","1000000001000000","1000000011001010","1000000011101000","1000000010000111","1000000011100100","1000000001111010","1000000001100010","1000000011011001","1000001001010000","1000000100000101","1000000000111100","0000000010010111","0000000010010111","1000000000001101","0000000101011010","1000000000010100","0000000000110110","0000000000101000","0000000000010101","0000000010010011","0000000001010111","0000000011010100","0000000011000010","0000000001101011","0000000001110101","0000000001010000","0000000010111101","0000000011100000","0000000000111011","1000000001000011","1000000000101110","1000000001001000","1000000000010110","1000000000000011","0000000000101101","1000000000010101","1000000101010001","1000000011111011","1000000000010101","0000000010111001","0000000000100110","1000000001101011","0000000101101010","0000000010001110","0000000100101101","0000000001011000","0000000011101110","0000000001110011","0000000001111001","0000000011001101","0000000001010100","0000000001101011","0000000000010100","0000000000101010","0000000010100010","0000000100010111","0000000010010101","0000000001000110","1000000000000111","1000000001011110","0000000000000010","0000000001001001","0000000010111110","0000000100001111","1000000000110000","1000000000010101","1000000010101010","1000000000011011","0000000001100010","1000000010010000","0000000000001101","0000000000111111","0000000011010111","0000000011011101","0000000100000110","0000000001100110","0000000001010100","0000000000111001","0000000000011100","1000000001011010","1000000001010001","0000000001010110","0000000011000011","0000000100100100","0000000011000100","0000000000100001","1000000000000000","0000000000000100","0000000000101100","0000000000101010","0000000001001011","0000000001100000","0000000001111010","0000000000101101","1000000101010100","1000000010110100","0000000001101101","0000000010110001","0000000001100111","0000000001010010","0000000010011100","0000000010110000","0000000001011101","0000000010000010","0000000011000001","0000000001110101","1000000000010111","1000000001111110","1000000000010000","0000000001011100","0000000011001000","0000000011111111","0000000010110001","0000000000100111","1000000000010000","0000000000011101","0000000000111100","0000000001111100","0000000011011000","0000000001010010","0000000000111110","0000000010010011","1000000100100101","1000000010111011","0000000010110010","0000000000001110","0000000001010101","1000000010110000","1000000011110010","1000000010000000","0000000000000100","0000000011000110","0000000010000101","0000000001011000","0000000000000000","0000000001111000","0000000000010100","0000000001011110","0000000011111000","0000000010001001","0000000010101010","0000000000110001","1000000000100001","0000000000100001","0000000001101110","0000000001011011","0000000010100001","0000000001111011","1000000000010001","1000000001111011","1000000011010011","1000000001010001","0000000010000001","0000000010000001","0000000001100010","1000000101100000","1000000100101101","1000000100011010","1000000000000000","0000000010000011","0000000010011010","0000000001011100","0000000010000001","0000000010010011","1000000000100101","0000000001110010","0000000100011110","0000000001110001","0000000000110000","1000000010000101","1000000001000011","0000000000100001","0000000000100111","0000000000001001","0000000000100101","0000000000010010","1000000001100011","1000000001001111","1000000010000111","1000000001001010","0000000000010001","0000000001110100","0000000010011001","1000000101010000","1000000101000010","1000000011100111","1000000001010110","1000000000001111","0000000001010101","0000000001110110","0000000100000000","0000000010000111","0000000001001000","0000000011110001","0000000101001101","0000000010001001","1000000000101010","1000000001110100","1000000001100001","1000000001110010","1000000001101100","1000000000100010","1000000000011111","1000000010001010","1000000011000001","0000000010110010","1000000010010001","1000000011001101","1000000000001111","0000000001101011","0000000011110010","1000000001111000","1000000100101010","1000000101100111","1000000010111011","1000000010000101","0000000000010110","0000000000100111","0000000000110001","0000000001001111","0000000001010001","0000000001111101","0000000011001100","0000000001010011","1000000001000000","1000000010001000","1000000000011110","1000000000110100","0000000000010011","1000000001001110","1000000001111110","1000000011010010","1000000100001010","0000000001010011","0000000010011111","0000000001100000","0000000001110101","1000000010001101","1000000000110111","1000000001100010","1000000010000100","1000000101000011","1000000010111001","1000000001011000","1000000010010110","1000000001010001","1000000001100111","0000000000010000","1000000000000001","0000000001111101","0000000001011100","0000000000001010","0000000000011010","1000000000101100","1000000001010111","0000000000100100","0000000001100010","1000000000001011","1000000010111111","1000000011010011","1000000010011000","1000000001010101","0000000000110011","0000000010100100","1000000000001111","1000000010011010","1000000001101010","1000000110010010","1000000010101010","1000000010101010","1000000010000110","1000000010110100","1000000001011011","1000000001001110","1000000001110001","1000000000110101","1000000000010110","0000000001000010","0000000010101101","0000000000011000","0000000010000000","0000000001000101","0000000000011001","1000000000001001","1000000000111101","1000000000011101","1000000001111111","1000000010010111","1000000000011110","0000000000000000","0000000000111010","0000000001000000","0000000010001010","0000000000010110","1000000010000100","1000000011000010","1000000011111011","1000000001010101","1000000010110110","1000000001111110","1000000001101111","1000000000010111","1000000000000010","1000000000110001","1000000000101000","0000000000101101","0000000001000010","1000000000001110","1000000000000111","0000000000001011","1000000001001011","1000000000011100","0000000000101000","1000000000001000","1000000000110000","1000000010100100","0000000001111001","0000000000010100","1000000001110111","1000000000001010","0000000001100000","0000000001101001","0000000000111010","1000000001101110","1000000000011111","1000000000010100","1000000001100100","1000000001010001","1000000001110001","1000000000111100","1000000001001100","1000000010100111","1000000001100000","1000000001101010","1000000000001000","0000000000000100","1000000000001010","0000000000000010","1000000000010111","0000000000101100","0000000000110010","0000000000000001","1000000010111101","1000000000100110","0000000001001010","0000000000110100","0000000001101011","1000000000110000","1000000000001000","1000000000010011","1000000000011001","1000000001111000","1000000000000100","0000000000100110","1000000000100110","1000000001110110","1000000000111101","1000000000000000","1000000010110001","1000000011110001","1000000001011100","1000000010010111","1000000001111111","1000000000101000","1000000000001010","1000000000010000","0000000000001100","0000000000000010","0000000000100000","1000000000110100","1000000001011011","1000000001010100","1000000000010111","1000000100001101","0000000010010100","1000000000010010","0000000000010011","1000000000000011","1000000010100011","1000000100000111","0000000001001010","1000000000101101","1000000001010110","1000000000101100","1000000000111100","0000000000110011","1000000001000000","1000000010011110","1000000011101101","1000000100011111","1000000100011010","1000000011110011","1000000011000111","1000000001110000","0000000000001110","1000000000001110","0000000001100000","0000000001010110","1000000000000000","0000000010111100","1000000000111101","1000000000110011","0000000000000110","1000000000001010","0000000000010110","1000000000001000","0000000001110100","0000000011001000","0000000000111100","0000000000001001","1000000010000100","1000000000011000","1000000000010110","1000000000100110","1000000010001011","1000000011001101","1000000001011001","0000000000010111","0000000010110111","0000000000000100","1000000100001110","1000000100010111","1000000010011000","1000000010011011","1000000001000000","1000000000011010","1000000001010011","1000000010010111","0000000000111111","1000000001100001","1000000010000101","0000000000001100","0000000000010011","0000000000000011","0000000000001010","0000000001101011","0000000011000001","0000000100001110","0000000111001110","0000000010111010","0000000010011101","0000000011111011","0000000010011101","0000000010001100","0000000001101101","0000000010011100","0000000100101100","0000000001010011","1000000001111000","1000000000101110","1000000001001010","1000000001110000","1000000001011100","0000000000010010","1000000001000001","0000000001011001","0000000000000001","0000000001110001","0000000000000111","0000000000000001","1000000000001100","1000000000010001","0000000000010001","1000000000000000","1000000000010000","0000000000110100","0000000011000010","0000000010101011","0000000100001111","0000000101000100","0000000010101010","0000000010100010","0000000001001000","0000000010100111","0000000101110110","0000000101100110","0000000010100111","0000000000100010","0000000010010111","0000000000111001","0000000001001111","0000000001011101","0000000001110001","1000000001111000","1000000000010010","1000000000001011","0000000000010010","1000000000010000");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
