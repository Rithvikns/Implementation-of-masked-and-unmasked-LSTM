library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity fully_connected_layer_0 is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_0 : out STD_LOGIC_VECTOR(15 downto 0);
        y_1 : out STD_LOGIC_VECTOR(15 downto 0);
        y_2 : out STD_LOGIC_VECTOR(15 downto 0);
        y_3 : out STD_LOGIC_VECTOR(15 downto 0);
        y_4 : out STD_LOGIC_VECTOR(15 downto 0);
        y_5 : out STD_LOGIC_VECTOR(15 downto 0);
        y_6 : out STD_LOGIC_VECTOR(15 downto 0);
        y_7 : out STD_LOGIC_VECTOR(15 downto 0);
        y_8 : out STD_LOGIC_VECTOR(15 downto 0);
        y_9 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end fully_connected_layer_0 ;
architecture Behavioral of fully_connected_layer_0 is

component fully_connected_layer_0_0  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_0 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_1  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_1 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_2  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_2 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_3  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_3 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_4  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_4 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_5  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_5 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_6  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_6 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_7  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_7 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_8  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_8 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;
component fully_connected_layer_0_9  is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_9 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component ;


 
begin
ut0_fully_connected_layer_0_0: fully_connected_layer_0_0 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_0 => y_0 
    );
ut1_fully_connected_layer_0_1: fully_connected_layer_0_1 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_1 => y_1 
    );
ut2_fully_connected_layer_0_2: fully_connected_layer_0_2 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_2 => y_2 
    );
ut3_fully_connected_layer_0_3: fully_connected_layer_0_3 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_3 => y_3 
    );
ut4_fully_connected_layer_0_4: fully_connected_layer_0_4 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_4 => y_4 
    );
ut5_fully_connected_layer_0_5: fully_connected_layer_0_5 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_5 => y_5 
    );
ut6_fully_connected_layer_0_6: fully_connected_layer_0_6 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_6 => y_6 
    );
ut7_fully_connected_layer_0_7: fully_connected_layer_0_7 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_7 => y_7 
    );
ut8_fully_connected_layer_0_8: fully_connected_layer_0_8 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_8 => y_8 
    );
ut9_fully_connected_layer_0_9: fully_connected_layer_0_9 port map(
clk => clk,
x_0 => x_0 ,
x_1 => x_1 ,
x_2 => x_2 ,
x_3 => x_3 ,
x_4 => x_4 ,
x_5 => x_5 ,
x_6 => x_6 ,
x_7 => x_7 ,
x_8 => x_8 ,
x_9 => x_9 ,
x_10 => x_10 ,
x_11 => x_11 ,
x_12 => x_12 ,
x_13 => x_13 ,
x_14 => x_14 ,
x_15 => x_15 ,
x_16 => x_16 ,
x_17 => x_17 ,
x_18 => x_18 ,
x_19 => x_19 ,
x_20 => x_20 ,
x_21 => x_21 ,
x_22 => x_22 ,
x_23 => x_23 ,
x_24 => x_24 ,
x_25 => x_25 ,
x_26 => x_26 ,
x_27 => x_27 ,
x_28 => x_28 ,
x_29 => x_29 ,
x_30 => x_30 ,
x_31 => x_31 ,
x_32 => x_32 ,
x_33 => x_33 ,
x_34 => x_34 ,
x_35 => x_35 ,
x_36 => x_36 ,
x_37 => x_37 ,
x_38 => x_38 ,
x_39 => x_39 ,
x_40 => x_40 ,
x_41 => x_41 ,
x_42 => x_42 ,
x_43 => x_43 ,
x_44 => x_44 ,
x_45 => x_45 ,
x_46 => x_46 ,
x_47 => x_47 ,
x_48 => x_48 ,
x_49 => x_49 ,
x_50 => x_50 ,
x_51 => x_51 ,
x_52 => x_52 ,
x_53 => x_53 ,
x_54 => x_54 ,
x_55 => x_55 ,
x_56 => x_56 ,
x_57 => x_57 ,
x_58 => x_58 ,
x_59 => x_59 ,
x_60 => x_60 ,
x_61 => x_61 ,
x_62 => x_62 ,
x_63 => x_63 ,
x_64 => x_64 ,
x_65 => x_65 ,
x_66 => x_66 ,
x_67 => x_67 ,
x_68 => x_68 ,
x_69 => x_69 ,
x_70 => x_70 ,
x_71 => x_71 ,
x_72 => x_72 ,
x_73 => x_73 ,
x_74 => x_74 ,
x_75 => x_75 ,
x_76 => x_76 ,
x_77 => x_77 ,
x_78 => x_78 ,
x_79 => x_79 ,
x_80 => x_80 ,
x_81 => x_81 ,
x_82 => x_82 ,
x_83 => x_83 ,
x_84 => x_84 ,
x_85 => x_85 ,
x_86 => x_86 ,
x_87 => x_87 ,
x_88 => x_88 ,
x_89 => x_89 ,
x_90 => x_90 ,
x_91 => x_91 ,
x_92 => x_92 ,
x_93 => x_93 ,
x_94 => x_94 ,
x_95 => x_95 ,
x_96 => x_96 ,
x_97 => x_97 ,
x_98 => x_98 ,
x_99 => x_99 ,
x_100 => x_100 ,
x_101 => x_101 ,
x_102 => x_102 ,
x_103 => x_103 ,
x_104 => x_104 ,
x_105 => x_105 ,
x_106 => x_106 ,
x_107 => x_107 ,
x_108 => x_108 ,
x_109 => x_109 ,
x_110 => x_110 ,
x_111 => x_111 ,
x_112 => x_112 ,
x_113 => x_113 ,
x_114 => x_114 ,
x_115 => x_115 ,
x_116 => x_116 ,
x_117 => x_117 ,
x_118 => x_118 ,
x_119 => x_119 ,
x_120 => x_120 ,
x_121 => x_121 ,
x_122 => x_122 ,
x_123 => x_123 ,
x_124 => x_124 ,
x_125 => x_125 ,
x_126 => x_126 ,
x_127 => x_127 ,
x_128 => x_128 ,
x_129 => x_129 ,
x_130 => x_130 ,
x_131 => x_131 ,
x_132 => x_132 ,
x_133 => x_133 ,
x_134 => x_134 ,
x_135 => x_135 ,
x_136 => x_136 ,
x_137 => x_137 ,
x_138 => x_138 ,
x_139 => x_139 ,
x_140 => x_140 ,
x_141 => x_141 ,
x_142 => x_142 ,
x_143 => x_143 ,
x_144 => x_144 ,
x_145 => x_145 ,
x_146 => x_146 ,
x_147 => x_147 ,
x_148 => x_148 ,
x_149 => x_149 ,
x_150 => x_150 ,
x_151 => x_151 ,
x_152 => x_152 ,
x_153 => x_153 ,
x_154 => x_154 ,
x_155 => x_155 ,
x_156 => x_156 ,
x_157 => x_157 ,
x_158 => x_158 ,
x_159 => x_159 ,
x_160 => x_160 ,
x_161 => x_161 ,
x_162 => x_162 ,
x_163 => x_163 ,
x_164 => x_164 ,
x_165 => x_165 ,
x_166 => x_166 ,
x_167 => x_167 ,
x_168 => x_168 ,
x_169 => x_169 ,
x_170 => x_170 ,
x_171 => x_171 ,
x_172 => x_172 ,
x_173 => x_173 ,
x_174 => x_174 ,
x_175 => x_175 ,
x_176 => x_176 ,
x_177 => x_177 ,
x_178 => x_178 ,
x_179 => x_179 ,
x_180 => x_180 ,
x_181 => x_181 ,
x_182 => x_182 ,
x_183 => x_183 ,
x_184 => x_184 ,
x_185 => x_185 ,
x_186 => x_186 ,
x_187 => x_187 ,
x_188 => x_188 ,
x_189 => x_189 ,
x_190 => x_190 ,
x_191 => x_191 ,
x_192 => x_192 ,
x_193 => x_193 ,
x_194 => x_194 ,
x_195 => x_195 ,
x_196 => x_196 ,
x_197 => x_197 ,
x_198 => x_198 ,
x_199 => x_199 ,
x_200 => x_200 ,
x_201 => x_201 ,
x_202 => x_202 ,
x_203 => x_203 ,
x_204 => x_204 ,
x_205 => x_205 ,
x_206 => x_206 ,
x_207 => x_207 ,
x_208 => x_208 ,
x_209 => x_209 ,
x_210 => x_210 ,
x_211 => x_211 ,
x_212 => x_212 ,
x_213 => x_213 ,
x_214 => x_214 ,
x_215 => x_215 ,
x_216 => x_216 ,
x_217 => x_217 ,
x_218 => x_218 ,
x_219 => x_219 ,
x_220 => x_220 ,
x_221 => x_221 ,
x_222 => x_222 ,
x_223 => x_223 ,
x_224 => x_224 ,
x_225 => x_225 ,
x_226 => x_226 ,
x_227 => x_227 ,
x_228 => x_228 ,
x_229 => x_229 ,
x_230 => x_230 ,
x_231 => x_231 ,
x_232 => x_232 ,
x_233 => x_233 ,
x_234 => x_234 ,
x_235 => x_235 ,
x_236 => x_236 ,
x_237 => x_237 ,
x_238 => x_238 ,
x_239 => x_239 ,
x_240 => x_240 ,
x_241 => x_241 ,
x_242 => x_242 ,
x_243 => x_243 ,
x_244 => x_244 ,
x_245 => x_245 ,
x_246 => x_246 ,
x_247 => x_247 ,
x_248 => x_248 ,
x_249 => x_249 ,
x_250 => x_250 ,
x_251 => x_251 ,
x_252 => x_252 ,
x_253 => x_253 ,
x_254 => x_254 ,
x_255 => x_255 ,
x_256 => x_256 ,
x_257 => x_257 ,
x_258 => x_258 ,
x_259 => x_259 ,
x_260 => x_260 ,
x_261 => x_261 ,
x_262 => x_262 ,
x_263 => x_263 ,
x_264 => x_264 ,
x_265 => x_265 ,
x_266 => x_266 ,
x_267 => x_267 ,
x_268 => x_268 ,
x_269 => x_269 ,
x_270 => x_270 ,
x_271 => x_271 ,
x_272 => x_272 ,
x_273 => x_273 ,
x_274 => x_274 ,
x_275 => x_275 ,
x_276 => x_276 ,
x_277 => x_277 ,
x_278 => x_278 ,
x_279 => x_279 ,
x_280 => x_280 ,
x_281 => x_281 ,
x_282 => x_282 ,
x_283 => x_283 ,
x_284 => x_284 ,
x_285 => x_285 ,
x_286 => x_286 ,
x_287 => x_287 ,
x_288 => x_288 ,
x_289 => x_289 ,
x_290 => x_290 ,
x_291 => x_291 ,
x_292 => x_292 ,
x_293 => x_293 ,
x_294 => x_294 ,
x_295 => x_295 ,
x_296 => x_296 ,
x_297 => x_297 ,
x_298 => x_298 ,
x_299 => x_299 ,
x_300 => x_300 ,
x_301 => x_301 ,
x_302 => x_302 ,
x_303 => x_303 ,
x_304 => x_304 ,
x_305 => x_305 ,
x_306 => x_306 ,
x_307 => x_307 ,
x_308 => x_308 ,
x_309 => x_309 ,
x_310 => x_310 ,
x_311 => x_311 ,
x_312 => x_312 ,
x_313 => x_313 ,
x_314 => x_314 ,
x_315 => x_315 ,
x_316 => x_316 ,
x_317 => x_317 ,
x_318 => x_318 ,
x_319 => x_319 ,
x_320 => x_320 ,
x_321 => x_321 ,
x_322 => x_322 ,
x_323 => x_323 ,
x_324 => x_324 ,
x_325 => x_325 ,
x_326 => x_326 ,
x_327 => x_327 ,
x_328 => x_328 ,
x_329 => x_329 ,
x_330 => x_330 ,
x_331 => x_331 ,
x_332 => x_332 ,
x_333 => x_333 ,
x_334 => x_334 ,
x_335 => x_335 ,
x_336 => x_336 ,
x_337 => x_337 ,
x_338 => x_338 ,
x_339 => x_339 ,
x_340 => x_340 ,
x_341 => x_341 ,
x_342 => x_342 ,
x_343 => x_343 ,
x_344 => x_344 ,
x_345 => x_345 ,
x_346 => x_346 ,
x_347 => x_347 ,
x_348 => x_348 ,
x_349 => x_349 ,
x_350 => x_350 ,
x_351 => x_351 ,
x_352 => x_352 ,
x_353 => x_353 ,
x_354 => x_354 ,
x_355 => x_355 ,
x_356 => x_356 ,
x_357 => x_357 ,
x_358 => x_358 ,
x_359 => x_359 ,
x_360 => x_360 ,
x_361 => x_361 ,
x_362 => x_362 ,
x_363 => x_363 ,
x_364 => x_364 ,
x_365 => x_365 ,
x_366 => x_366 ,
x_367 => x_367 ,
x_368 => x_368 ,
x_369 => x_369 ,
x_370 => x_370 ,
x_371 => x_371 ,
x_372 => x_372 ,
x_373 => x_373 ,
x_374 => x_374 ,
x_375 => x_375 ,
x_376 => x_376 ,
x_377 => x_377 ,
x_378 => x_378 ,
x_379 => x_379 ,
x_380 => x_380 ,
x_381 => x_381 ,
x_382 => x_382 ,
x_383 => x_383 ,
x_384 => x_384 ,
x_385 => x_385 ,
x_386 => x_386 ,
x_387 => x_387 ,
x_388 => x_388 ,
x_389 => x_389 ,
x_390 => x_390 ,
x_391 => x_391 ,
x_392 => x_392 ,
x_393 => x_393 ,
x_394 => x_394 ,
x_395 => x_395 ,
x_396 => x_396 ,
x_397 => x_397 ,
x_398 => x_398 ,
x_399 => x_399 ,
x_400 => x_400 ,
x_401 => x_401 ,
x_402 => x_402 ,
x_403 => x_403 ,
x_404 => x_404 ,
x_405 => x_405 ,
x_406 => x_406 ,
x_407 => x_407 ,
x_408 => x_408 ,
x_409 => x_409 ,
x_410 => x_410 ,
x_411 => x_411 ,
x_412 => x_412 ,
x_413 => x_413 ,
x_414 => x_414 ,
x_415 => x_415 ,
x_416 => x_416 ,
x_417 => x_417 ,
x_418 => x_418 ,
x_419 => x_419 ,
x_420 => x_420 ,
x_421 => x_421 ,
x_422 => x_422 ,
x_423 => x_423 ,
x_424 => x_424 ,
x_425 => x_425 ,
x_426 => x_426 ,
x_427 => x_427 ,
x_428 => x_428 ,
x_429 => x_429 ,
x_430 => x_430 ,
x_431 => x_431 ,
x_432 => x_432 ,
x_433 => x_433 ,
x_434 => x_434 ,
x_435 => x_435 ,
x_436 => x_436 ,
x_437 => x_437 ,
x_438 => x_438 ,
x_439 => x_439 ,
x_440 => x_440 ,
x_441 => x_441 ,
x_442 => x_442 ,
x_443 => x_443 ,
x_444 => x_444 ,
x_445 => x_445 ,
x_446 => x_446 ,
x_447 => x_447 ,
x_448 => x_448 ,
x_449 => x_449 ,
x_450 => x_450 ,
x_451 => x_451 ,
x_452 => x_452 ,
x_453 => x_453 ,
x_454 => x_454 ,
x_455 => x_455 ,
x_456 => x_456 ,
x_457 => x_457 ,
x_458 => x_458 ,
x_459 => x_459 ,
x_460 => x_460 ,
x_461 => x_461 ,
x_462 => x_462 ,
x_463 => x_463 ,
x_464 => x_464 ,
x_465 => x_465 ,
x_466 => x_466 ,
x_467 => x_467 ,
x_468 => x_468 ,
x_469 => x_469 ,
x_470 => x_470 ,
x_471 => x_471 ,
x_472 => x_472 ,
x_473 => x_473 ,
x_474 => x_474 ,
x_475 => x_475 ,
x_476 => x_476 ,
x_477 => x_477 ,
x_478 => x_478 ,
x_479 => x_479 ,
x_480 => x_480 ,
x_481 => x_481 ,
x_482 => x_482 ,
x_483 => x_483 ,
x_484 => x_484 ,
x_485 => x_485 ,
x_486 => x_486 ,
x_487 => x_487 ,
x_488 => x_488 ,
x_489 => x_489 ,
x_490 => x_490 ,
x_491 => x_491 ,
x_492 => x_492 ,
x_493 => x_493 ,
x_494 => x_494 ,
x_495 => x_495 ,
x_496 => x_496 ,
x_497 => x_497 ,
x_498 => x_498 ,
x_499 => x_499 ,
x_500 => x_500 ,
x_501 => x_501 ,
x_502 => x_502 ,
x_503 => x_503 ,
x_504 => x_504 ,
x_505 => x_505 ,
x_506 => x_506 ,
x_507 => x_507 ,
x_508 => x_508 ,
x_509 => x_509 ,
x_510 => x_510 ,
x_511 => x_511 ,
x_512 => x_512 ,
x_513 => x_513 ,
x_514 => x_514 ,
x_515 => x_515 ,
x_516 => x_516 ,
x_517 => x_517 ,
x_518 => x_518 ,
x_519 => x_519 ,
x_520 => x_520 ,
x_521 => x_521 ,
x_522 => x_522 ,
x_523 => x_523 ,
x_524 => x_524 ,
x_525 => x_525 ,
x_526 => x_526 ,
x_527 => x_527 ,
x_528 => x_528 ,
x_529 => x_529 ,
x_530 => x_530 ,
x_531 => x_531 ,
x_532 => x_532 ,
x_533 => x_533 ,
x_534 => x_534 ,
x_535 => x_535 ,
x_536 => x_536 ,
x_537 => x_537 ,
x_538 => x_538 ,
x_539 => x_539 ,
x_540 => x_540 ,
x_541 => x_541 ,
x_542 => x_542 ,
x_543 => x_543 ,
x_544 => x_544 ,
x_545 => x_545 ,
x_546 => x_546 ,
x_547 => x_547 ,
x_548 => x_548 ,
x_549 => x_549 ,
x_550 => x_550 ,
x_551 => x_551 ,
x_552 => x_552 ,
x_553 => x_553 ,
x_554 => x_554 ,
x_555 => x_555 ,
x_556 => x_556 ,
x_557 => x_557 ,
x_558 => x_558 ,
x_559 => x_559 ,
x_560 => x_560 ,
x_561 => x_561 ,
x_562 => x_562 ,
x_563 => x_563 ,
x_564 => x_564 ,
x_565 => x_565 ,
x_566 => x_566 ,
x_567 => x_567 ,
x_568 => x_568 ,
x_569 => x_569 ,
x_570 => x_570 ,
x_571 => x_571 ,
x_572 => x_572 ,
x_573 => x_573 ,
x_574 => x_574 ,
x_575 => x_575 ,
x_576 => x_576 ,
x_577 => x_577 ,
x_578 => x_578 ,
x_579 => x_579 ,
x_580 => x_580 ,
x_581 => x_581 ,
x_582 => x_582 ,
x_583 => x_583 ,
x_584 => x_584 ,
x_585 => x_585 ,
x_586 => x_586 ,
x_587 => x_587 ,
x_588 => x_588 ,
x_589 => x_589 ,
x_590 => x_590 ,
x_591 => x_591 ,
x_592 => x_592 ,
x_593 => x_593 ,
x_594 => x_594 ,
x_595 => x_595 ,
x_596 => x_596 ,
x_597 => x_597 ,
x_598 => x_598 ,
x_599 => x_599 ,
x_600 => x_600 ,
x_601 => x_601 ,
x_602 => x_602 ,
x_603 => x_603 ,
x_604 => x_604 ,
x_605 => x_605 ,
x_606 => x_606 ,
x_607 => x_607 ,
x_608 => x_608 ,
x_609 => x_609 ,
x_610 => x_610 ,
x_611 => x_611 ,
x_612 => x_612 ,
x_613 => x_613 ,
x_614 => x_614 ,
x_615 => x_615 ,
x_616 => x_616 ,
x_617 => x_617 ,
x_618 => x_618 ,
x_619 => x_619 ,
x_620 => x_620 ,
x_621 => x_621 ,
x_622 => x_622 ,
x_623 => x_623 ,
x_624 => x_624 ,
x_625 => x_625 ,
x_626 => x_626 ,
x_627 => x_627 ,
x_628 => x_628 ,
x_629 => x_629 ,
x_630 => x_630 ,
x_631 => x_631 ,
x_632 => x_632 ,
x_633 => x_633 ,
x_634 => x_634 ,
x_635 => x_635 ,
x_636 => x_636 ,
x_637 => x_637 ,
x_638 => x_638 ,
x_639 => x_639 ,
x_640 => x_640 ,
x_641 => x_641 ,
x_642 => x_642 ,
x_643 => x_643 ,
x_644 => x_644 ,
x_645 => x_645 ,
x_646 => x_646 ,
x_647 => x_647 ,
x_648 => x_648 ,
x_649 => x_649 ,
x_650 => x_650 ,
x_651 => x_651 ,
x_652 => x_652 ,
x_653 => x_653 ,
x_654 => x_654 ,
x_655 => x_655 ,
x_656 => x_656 ,
x_657 => x_657 ,
x_658 => x_658 ,
x_659 => x_659 ,
x_660 => x_660 ,
x_661 => x_661 ,
x_662 => x_662 ,
x_663 => x_663 ,
x_664 => x_664 ,
x_665 => x_665 ,
x_666 => x_666 ,
x_667 => x_667 ,
x_668 => x_668 ,
x_669 => x_669 ,
x_670 => x_670 ,
x_671 => x_671 ,
x_672 => x_672 ,
x_673 => x_673 ,
x_674 => x_674 ,
x_675 => x_675 ,
x_676 => x_676 ,
x_677 => x_677 ,
x_678 => x_678 ,
x_679 => x_679 ,
x_680 => x_680 ,
x_681 => x_681 ,
x_682 => x_682 ,
x_683 => x_683 ,
x_684 => x_684 ,
x_685 => x_685 ,
x_686 => x_686 ,
x_687 => x_687 ,
x_688 => x_688 ,
x_689 => x_689 ,
x_690 => x_690 ,
x_691 => x_691 ,
x_692 => x_692 ,
x_693 => x_693 ,
x_694 => x_694 ,
x_695 => x_695 ,
x_696 => x_696 ,
x_697 => x_697 ,
x_698 => x_698 ,
x_699 => x_699 ,
x_700 => x_700 ,
x_701 => x_701 ,
x_702 => x_702 ,
x_703 => x_703 ,
x_704 => x_704 ,
x_705 => x_705 ,
x_706 => x_706 ,
x_707 => x_707 ,
x_708 => x_708 ,
x_709 => x_709 ,
x_710 => x_710 ,
x_711 => x_711 ,
x_712 => x_712 ,
x_713 => x_713 ,
x_714 => x_714 ,
x_715 => x_715 ,
x_716 => x_716 ,
x_717 => x_717 ,
x_718 => x_718 ,
x_719 => x_719 ,
x_720 => x_720 ,
x_721 => x_721 ,
x_722 => x_722 ,
x_723 => x_723 ,
x_724 => x_724 ,
x_725 => x_725 ,
x_726 => x_726 ,
x_727 => x_727 ,
x_728 => x_728 ,
x_729 => x_729 ,
x_730 => x_730 ,
x_731 => x_731 ,
x_732 => x_732 ,
x_733 => x_733 ,
x_734 => x_734 ,
x_735 => x_735 ,
x_736 => x_736 ,
x_737 => x_737 ,
x_738 => x_738 ,
x_739 => x_739 ,
x_740 => x_740 ,
x_741 => x_741 ,
x_742 => x_742 ,
x_743 => x_743 ,
x_744 => x_744 ,
x_745 => x_745 ,
x_746 => x_746 ,
x_747 => x_747 ,
x_748 => x_748 ,
x_749 => x_749 ,
x_750 => x_750 ,
x_751 => x_751 ,
x_752 => x_752 ,
x_753 => x_753 ,
x_754 => x_754 ,
x_755 => x_755 ,
x_756 => x_756 ,
x_757 => x_757 ,
x_758 => x_758 ,
x_759 => x_759 ,
x_760 => x_760 ,
x_761 => x_761 ,
x_762 => x_762 ,
x_763 => x_763 ,
x_764 => x_764 ,
x_765 => x_765 ,
x_766 => x_766 ,
x_767 => x_767 ,
x_768 => x_768 ,
x_769 => x_769 ,
x_770 => x_770 ,
x_771 => x_771 ,
x_772 => x_772 ,
x_773 => x_773 ,
x_774 => x_774 ,
x_775 => x_775 ,
x_776 => x_776 ,
x_777 => x_777 ,
x_778 => x_778 ,
x_779 => x_779 ,
x_780 => x_780 ,
x_781 => x_781 ,
x_782 => x_782 ,
x_783 => x_783 ,
y_9 => y_9 
    );

end Behavioral;