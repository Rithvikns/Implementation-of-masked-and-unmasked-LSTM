library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity raminfr is
port (
        clk : in std_logic;
        we : in std_logic;
        a : in std_logic_vector(8 downto 0);
        di : in std_logic_vector(7 downto 0);
        do : out std_logic_vector(7 downto 0)
    );
end raminfr;

architecture syn of raminfr is

type ram_type is array (0 to 489) of std_logic_vector (7 downto 0);


signal RAM : ram_type := ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11011000","10011011","11111101","11111110","11111110","11010001","10110010","11100000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10001000","10110110","11111011","11111101","11111100","11111000","11111101","11111101","11111101","11101000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11000010","11111101","11110011","11100010","10010000","10010100","10110010","10110001","11111101","11101011","10011000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10010000","11110001","11111101","11110000","00000000","00000000","00000000","00000000","10011000","10111011","11111101","10100000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10001111","11111101","11000011","10100000","00000000","00000000","00000000","10010000","11100010","11111101","11111101","10101101","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10101110","11111101","10011110","00000000","00000000","00000000","00000000","10010000","11111101","11111101","11111101","11110110","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10000000","11001110","11111101","10001010","00000000","00000000","00000000","10000000","11100100","11111101","11111101","11110101","11001000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10101110","11111101","10001010","00000000","00000000","10000000","10100010","11111101","11111101","11000111","10000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10001001","11111101","10110001","10101100","00000000","10100100","11111101","11111101","11111101","11110100","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111000","11011100","11111101","11111011","11111001","11111101","11111101","11101011","11111101","10110111","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11010000","11000010","11111000","11111000","10111101","11010110","10011111","11111101","10110111","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10011111","11111101","10110111","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10011111","11111101","10111100","10000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10011111","11111101","11111101","11101000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10010000","11111101","11111101","11110000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11110000","11111101","11111101","10001010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
begin
process (clk)
    begin
    if (clk'event and clk = '1') then
    if (we = '1') then
    RAM(conv_integer(a)) <= di;
    end if;
    end if;
end process;
do <= RAM(conv_integer(a));
end syn;