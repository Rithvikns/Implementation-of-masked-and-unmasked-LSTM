library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity fully_connected_layer_1_7 is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        y_7 : out STD_LOGIC_VECTOR(15 downto 0)
    );
end fully_connected_layer_1_7 ;
architecture Behavioral of fully_connected_layer_1_7 is
signal store_sum : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_0 : STD_LOGIC_VECTOR(15 downto 0) := "1000001000000010";
signal store_weight_0 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_1 : STD_LOGIC_VECTOR(15 downto 0) := "0000001001000100";
signal store_weight_1 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_2 : STD_LOGIC_VECTOR(15 downto 0) := "1000000101110001";
signal store_weight_2 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_3 : STD_LOGIC_VECTOR(15 downto 0) := "1000011001110111";
signal store_weight_3 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_4 : STD_LOGIC_VECTOR(15 downto 0) := "1000010001000111";
signal store_weight_4 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_5 : STD_LOGIC_VECTOR(15 downto 0) := "0000000011100110";
signal store_weight_5 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_6 : STD_LOGIC_VECTOR(15 downto 0) := "0000001011100010";
signal store_weight_6 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_7 : STD_LOGIC_VECTOR(15 downto 0) := "1000010000000000";
signal store_weight_7 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_8 : STD_LOGIC_VECTOR(15 downto 0) := "1000000100101010";
signal store_weight_8 : STD_LOGIC_VECTOR(15 downto 0) ;
signal weight_9 : STD_LOGIC_VECTOR(15 downto 0) := "1000001101010000";
signal store_weight_9 : STD_LOGIC_VECTOR(15 downto 0) ;
signal sum_0 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_1 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_2 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_3 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_4 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_5 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_6 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_7 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_8 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_9 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_10 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_11 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_12 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_13 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_14 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_15 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_16 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_17 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_18 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_19 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_20 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_21 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_22 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_23 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_24 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_25 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_26 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_27 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_28 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_29 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_30 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_31 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_32 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_33 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_34 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_35 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_36 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_37 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_38 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_39 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_40 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_41 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_42 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_43 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_44 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_45 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_46 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_47 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_48 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_49 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_50 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_51 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_52 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_53 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_54 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_55 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_56 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_57 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_58 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_59 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_60 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_61 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_62 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_63 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_64 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_65 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_66 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_67 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_68 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_69 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_70 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_71 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_72 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_73 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_74 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_75 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_76 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_77 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_78 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_79 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_80 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_81 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_82 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_83 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_84 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_85 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_86 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_87 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_88 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_89 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_90 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_91 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_92 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_93 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_94 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_95 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_96 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_97 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_98 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_99 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_100 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_101 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_102 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_103 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_104 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_105 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_106 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_107 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_108 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_109 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_110 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_111 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_112 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_113 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_114 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_115 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_116 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_117 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_118 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_119 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_120 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_121 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_122 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_123 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_124 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_125 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_126 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_127 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_128 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_129 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_130 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_131 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_132 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_133 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_134 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_135 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_136 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_137 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_138 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_139 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_140 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_141 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_142 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_143 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_144 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_145 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_146 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_147 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_148 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_149 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_150 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_151 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_152 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_153 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_154 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_155 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_156 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_157 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_158 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_159 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_160 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_161 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_162 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_163 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_164 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_165 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_166 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_167 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_168 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_169 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_170 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_171 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_172 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_173 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_174 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_175 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_176 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_177 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_178 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_179 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_180 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_181 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_182 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_183 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_184 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_185 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_186 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_187 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_188 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_189 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_190 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_191 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_192 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_193 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_194 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_195 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_196 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_197 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_198 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_199 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_200 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_201 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_202 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_203 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_204 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_205 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_206 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_207 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_208 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_209 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_210 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_211 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_212 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_213 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_214 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_215 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_216 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_217 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_218 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_219 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_220 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_221 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_222 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_223 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_224 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_225 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_226 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_227 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_228 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_229 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_230 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_231 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_232 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_233 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_234 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_235 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_236 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_237 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_238 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_239 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_240 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_241 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_242 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_243 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_244 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_245 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_246 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_247 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_248 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_249 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_250 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_251 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_252 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_253 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_254 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_255 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_256 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_257 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_258 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_259 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_260 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_261 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_262 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_263 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_264 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_265 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_266 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_267 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_268 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_269 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_270 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_271 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_272 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_273 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_274 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_275 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_276 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_277 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_278 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_279 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_280 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_281 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_282 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_283 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_284 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_285 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_286 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_287 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_288 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_289 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_290 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_291 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_292 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_293 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_294 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_295 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_296 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_297 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_298 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_299 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_300 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_301 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_302 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_303 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_304 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_305 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_306 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_307 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_308 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_309 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_310 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_311 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_312 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_313 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_314 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_315 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_316 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_317 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_318 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_319 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_320 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_321 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_322 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_323 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_324 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_325 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_326 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_327 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_328 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_329 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_330 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_331 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_332 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_333 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_334 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_335 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_336 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_337 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_338 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_339 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_340 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_341 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_342 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_343 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_344 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_345 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_346 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_347 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_348 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_349 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_350 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_351 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_352 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_353 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_354 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_355 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_356 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_357 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_358 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_359 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_360 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_361 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_362 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_363 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_364 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_365 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_366 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_367 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_368 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_369 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_370 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_371 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_372 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_373 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_374 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_375 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_376 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_377 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_378 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_379 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_380 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_381 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_382 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_383 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_384 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_385 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_386 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_387 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_388 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_389 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_390 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_391 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_392 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_393 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_394 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_395 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_396 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_397 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_398 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_399 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_400 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_401 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_402 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_403 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_404 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_405 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_406 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_407 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_408 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_409 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_410 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_411 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_412 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_413 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_414 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_415 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_416 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_417 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_418 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_419 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_420 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_421 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_422 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_423 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_424 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_425 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_426 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_427 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_428 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_429 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_430 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_431 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_432 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_433 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_434 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_435 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_436 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_437 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_438 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_439 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_440 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_441 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_442 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_443 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_444 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_445 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_446 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_447 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_448 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_449 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_450 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_451 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_452 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_453 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_454 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_455 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_456 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_457 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_458 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_459 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_460 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_461 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_462 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_463 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_464 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_465 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_466 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_467 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_468 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_469 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_470 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_471 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_472 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_473 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_474 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_475 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_476 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_477 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_478 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_479 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_480 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_481 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_482 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_483 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_484 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_485 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_486 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_487 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_488 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_489 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_490 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_491 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_492 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_493 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_494 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_495 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_496 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_497 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_498 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_499 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_500 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_501 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_502 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_503 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_504 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_505 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_506 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_507 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_508 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_509 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_510 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_511 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_512 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_513 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_514 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_515 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_516 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_517 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_518 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_519 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_520 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_521 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_522 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_523 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_524 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_525 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_526 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_527 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_528 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_529 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_530 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_531 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_532 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_533 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_534 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_535 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_536 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_537 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_538 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_539 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_540 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_541 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_542 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_543 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_544 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_545 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_546 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_547 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_548 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_549 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_550 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_551 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_552 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_553 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_554 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_555 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_556 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_557 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_558 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_559 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_560 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_561 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_562 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_563 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_564 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_565 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_566 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_567 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_568 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_569 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_570 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_571 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_572 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_573 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_574 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_575 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_576 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_577 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_578 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_579 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_580 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_581 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_582 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_583 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_584 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_585 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_586 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_587 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_588 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_589 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_590 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_591 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_592 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_593 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_594 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_595 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_596 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_597 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_598 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_599 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_600 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_601 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_602 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_603 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_604 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_605 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_606 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_607 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_608 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_609 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_610 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_611 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_612 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_613 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_614 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_615 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_616 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_617 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_618 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_619 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_620 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_621 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_622 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_623 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_624 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_625 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_626 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_627 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_628 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_629 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_630 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_631 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_632 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_633 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_634 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_635 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_636 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_637 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_638 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_639 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_640 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_641 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_642 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_643 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_644 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_645 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_646 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_647 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_648 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_649 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_650 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_651 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_652 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_653 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_654 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_655 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_656 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_657 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_658 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_659 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_660 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_661 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_662 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_663 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_664 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_665 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_666 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_667 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_668 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_669 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_670 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_671 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_672 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_673 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_674 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_675 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_676 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_677 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_678 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_679 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_680 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_681 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_682 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_683 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_684 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_685 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_686 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_687 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_688 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_689 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_690 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_691 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_692 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_693 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_694 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_695 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_696 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_697 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_698 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_699 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_700 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_701 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_702 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_703 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_704 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_705 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_706 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_707 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_708 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_709 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_710 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_711 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_712 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_713 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_714 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_715 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_716 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_717 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_718 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_719 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_720 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_721 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_722 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_723 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_724 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_725 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_726 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_727 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_728 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_729 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_730 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_731 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_732 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_733 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_734 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_735 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_736 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_737 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_738 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_739 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_740 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_741 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_742 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_743 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_744 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_745 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_746 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_747 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_748 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_749 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_750 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_751 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_752 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_753 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_754 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_755 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_756 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_757 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_758 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_759 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_760 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_761 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_762 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_763 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_764 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_765 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_766 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_767 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_768 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_769 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_770 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_771 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_772 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_773 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_774 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_775 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_776 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_777 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_778 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_779 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_780 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_781 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal sum_782 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
signal biases : STD_LOGIC_VECTOR(15 downto 0) := "1000000100010011";
component  sigmoid is
	port (
		num:in integer ;
		y: out STD_LOGIC_VECTOR(15 downto 0)
		);
end component sigmoid;

component  nn_addition is
	Port (
		inputx : in STD_LOGIC_VECTOR(15 downto 0);
		inputy : in STD_LOGIC_VECTOR(15 downto 0);
		output : out STD_LOGIC_VECTOR(15 downto 0));
end component nn_addition;

component  nn_multiplication is
	Port (
		inputx : in STD_LOGIC_VECTOR(15 downto 0);
		inputy : in STD_LOGIC_VECTOR(15 downto 0);
		output : out STD_LOGIC_VECTOR(15 downto 0));
end component nn_multiplication;
begin
ut0_nn_multiplication: nn_multiplication port map(weight_0 , x_0 ,store_weight_0 );
ut1_nn_multiplication: nn_multiplication port map(weight_1 , x_1 ,store_weight_1 );
ut2_nn_multiplication: nn_multiplication port map(weight_2 , x_2 ,store_weight_2 );
ut3_nn_multiplication: nn_multiplication port map(weight_3 , x_3 ,store_weight_3 );
ut4_nn_multiplication: nn_multiplication port map(weight_4 , x_4 ,store_weight_4 );
ut5_nn_multiplication: nn_multiplication port map(weight_5 , x_5 ,store_weight_5 );
ut6_nn_multiplication: nn_multiplication port map(weight_6 , x_6 ,store_weight_6 );
ut7_nn_multiplication: nn_multiplication port map(weight_7 , x_7 ,store_weight_7 );
ut8_nn_multiplication: nn_multiplication port map(weight_8 , x_8 ,store_weight_8 );
ut9_nn_multiplication: nn_multiplication port map(weight_9 , x_9 ,store_weight_9 );
ut0_nn_addition: nn_addition port map( store_weight_0,store_weight_1,sum_0);
ut1_nn_addition: nn_addition port map( store_weight_2,store_weight_3,sum_1);
ut2_nn_addition: nn_addition port map( store_weight_4,store_weight_5,sum_2);
ut3_nn_addition: nn_addition port map( store_weight_6,store_weight_7,sum_3);
ut4_nn_addition: nn_addition port map( store_weight_8,store_weight_9,sum_4);
ut5_nn_addition: nn_addition port map( sum_0,sum_1,sum_5);
ut6_nn_addition: nn_addition port map( sum_2,sum_3,sum_6);
ut7_nn_addition: nn_addition port map( sum_4,sum_5,sum_7);
ut8_nn_addition: nn_addition port map( sum_6,sum_7,sum_8);
ut10_nn_addition: nn_addition port map(biases,sum_8 ,store_value);
ut1_sigmoid: sigmoid port map( to_integer(unsigned(store_value)),y_7);
end Behavioral;