library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity lstm is
    port (
        clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y : out STD_LOGIC_VECTOR(3 downto 0)
    );
end lstm ;

architecture Behavioral of lstm is

signal store_value_0 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_1 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_2 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_3 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_4 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_5 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_6 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_7 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_8 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_9 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_10 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_11 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_12 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_13 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_14 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_15 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_16 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_17 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_18 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_19 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_20 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_21 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_22 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_23 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_24 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_25 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_26 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_27 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_28 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_29 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_30 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_31 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_32 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_33 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_34 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_35 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_36 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_37 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_38 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_39 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_40 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_41 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_42 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_43 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_44 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_45 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_46 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_47 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_48 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_49 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_50 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_51 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_52 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_53 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_54 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_55 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_56 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_57 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_58 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_59 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_60 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_61 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_62 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_63 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_64 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_65 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_66 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_67 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_68 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_69 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_70 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_71 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_72 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_73 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_74 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_75 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_76 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_77 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_78 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_79 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_80 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_81 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_82 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_83 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_84 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_85 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_86 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_87 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_88 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_89 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_90 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_91 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_92 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_93 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_94 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_95 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_96 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_97 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_98 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_99 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_100 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_101 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_102 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_103 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_104 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_105 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_106 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_107 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_108 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_109 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_110 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_111 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_112 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_113 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_114 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_115 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_116 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_117 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_118 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_119 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_120 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_121 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_122 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_123 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_124 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_125 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_126 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_127 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_128 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_129 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_130 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_131 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_132 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_133 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_134 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_135 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_136 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_137 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_138 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_139 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_140 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_141 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_142 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_143 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_144 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_145 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_146 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_147 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_148 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_149 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_150 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_151 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_152 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_153 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_154 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_155 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_156 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_157 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_158 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_159 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_160 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_161 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_162 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_163 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_164 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_165 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_166 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_167 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_168 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_169 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_170 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_171 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_172 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_173 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_174 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_175 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_176 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_177 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_178 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_179 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_180 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_181 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_182 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_183 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_184 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_185 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_186 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_187 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_188 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_189 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_190 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_191 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_192 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_193 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_194 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_195 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_196 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_197 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_198 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_199 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_200 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_201 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_202 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_203 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_204 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_205 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_206 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_207 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_208 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_209 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_210 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_211 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_212 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_213 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_214 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_215 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_216 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_217 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_218 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_219 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_220 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_221 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_222 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_223 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_224 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_225 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_226 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_227 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_228 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_229 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_230 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_231 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_232 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_233 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_234 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_235 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_236 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_237 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_238 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_239 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_240 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_241 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_242 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_243 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_244 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_245 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_246 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_247 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_248 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_249 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_250 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_251 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_252 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_253 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_254 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_255 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_256 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_257 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_258 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_259 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_260 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_261 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_262 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_263 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_264 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_265 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_266 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_267 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_268 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_269 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_270 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_271 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_272 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_273 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_274 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_275 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_276 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_277 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_278 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_279 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_280 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_281 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_282 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_283 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_284 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_285 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_286 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_287 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_288 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_289 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_290 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_291 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_292 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_293 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_294 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_295 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_296 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_297 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_298 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_299 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_300 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_301 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_302 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_303 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_304 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_305 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_306 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_307 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_308 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_309 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_310 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_311 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_312 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_313 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_314 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_315 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_316 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_317 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_318 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_319 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_320 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_321 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_322 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_323 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_324 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_325 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_326 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_327 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_328 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_329 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_330 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_331 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_332 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_333 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_334 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_335 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_336 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_337 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_338 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_339 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_340 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_341 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_342 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_343 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_344 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_345 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_346 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_347 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_348 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_349 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_350 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_351 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_352 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_353 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_354 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_355 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_356 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_357 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_358 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_359 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_360 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_361 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_362 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_363 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_364 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_365 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_366 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_367 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_368 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_369 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_370 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_371 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_372 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_373 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_374 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_375 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_376 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_377 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_378 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_379 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_380 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_381 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_382 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_383 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_384 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_385 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_386 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_387 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_388 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_389 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_390 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_391 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_392 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_393 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_394 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_395 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_396 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_397 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_398 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_399 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_400 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_401 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_402 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_403 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_404 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_405 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_406 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_407 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_408 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_409 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_410 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_411 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_412 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_413 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_414 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_415 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_416 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_417 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_418 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_419 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_420 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_421 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_422 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_423 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_424 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_425 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_426 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_427 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_428 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_429 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_430 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_431 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_432 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_433 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_434 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_435 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_436 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_437 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_438 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_439 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_440 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_441 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_442 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_443 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_444 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_445 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_446 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_447 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_448 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_449 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_450 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_451 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_452 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_453 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_454 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_455 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_456 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_457 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_458 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_459 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_460 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_461 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_462 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_463 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_464 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_465 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_466 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_467 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_468 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_469 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_470 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_471 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_472 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_473 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_474 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_475 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_476 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_477 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_478 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_479 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_480 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_481 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_482 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_483 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_484 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_485 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_486 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_487 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_488 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_489 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_490 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_491 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_492 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_493 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_494 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_495 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_496 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_497 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_498 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_499 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_500 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_501 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_502 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_503 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_504 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_505 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_506 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_507 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_508 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_509 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_510 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_511 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_512 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_513 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_514 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_515 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_516 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_517 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_518 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_519 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_520 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_521 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_522 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_523 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_524 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_525 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_526 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_527 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_528 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_529 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_530 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_531 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_532 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_533 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_534 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_535 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_536 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_537 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_538 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_539 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_540 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_541 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_542 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_543 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_544 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_545 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_546 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_547 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_548 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_549 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_550 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_551 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_552 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_553 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_554 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_555 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_556 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_557 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_558 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_559 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_560 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_561 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_562 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_563 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_564 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_565 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_566 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_567 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_568 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_569 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_570 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_571 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_572 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_573 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_574 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_575 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_576 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_577 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_578 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_579 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_580 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_581 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_582 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_583 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_584 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_585 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_586 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_587 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_588 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_589 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_590 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_591 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_592 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_593 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_594 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_595 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_596 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_597 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_598 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_599 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_600 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_601 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_602 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_603 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_604 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_605 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_606 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_607 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_608 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_609 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_610 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_611 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_612 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_613 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_614 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_615 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_616 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_617 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_618 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_619 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_620 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_621 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_622 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_623 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_624 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_625 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_626 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_627 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_628 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_629 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_630 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_631 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_632 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_633 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_634 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_635 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_636 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_637 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_638 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_639 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_640 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_641 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_642 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_643 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_644 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_645 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_646 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_647 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_648 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_649 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_650 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_651 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_652 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_653 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_654 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_655 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_656 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_657 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_658 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_659 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_660 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_661 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_662 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_663 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_664 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_665 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_666 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_667 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_668 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_669 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_670 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_671 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_672 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_673 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_674 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_675 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_676 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_677 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_678 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_679 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_680 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_681 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_682 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_683 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_684 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_685 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_686 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_687 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_688 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_689 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_690 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_691 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_692 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_693 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_694 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_695 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_696 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_697 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_698 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_699 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_700 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_701 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_702 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_703 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_704 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_705 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_706 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_707 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_708 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_709 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_710 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_711 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_712 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_713 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_714 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_715 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_716 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_717 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_718 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_719 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_720 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_721 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_722 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_723 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_724 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_725 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_726 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_727 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_728 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_729 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_730 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_731 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_732 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_733 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_734 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_735 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_736 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_737 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_738 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_739 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_740 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_741 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_742 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_743 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_744 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_745 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_746 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_747 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_748 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_749 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_750 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_751 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_752 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_753 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_754 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_755 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_756 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_757 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_758 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_759 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_760 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_761 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_762 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_763 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_764 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_765 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_766 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_767 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_768 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_769 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_770 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_771 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_772 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_773 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_774 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_775 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_776 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_777 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_778 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_779 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_780 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_781 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_782 : STD_LOGIC_VECTOR(15 downto 0) ;
signal store_value_783 : STD_LOGIC_VECTOR(15 downto 0) ;

component  lstm_layer is
	Port (
		clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y_0 : out STD_LOGIC_VECTOR(15 downto 0);
        y_1 : out STD_LOGIC_VECTOR(15 downto 0);
        y_2 : out STD_LOGIC_VECTOR(15 downto 0);
        y_3 : out STD_LOGIC_VECTOR(15 downto 0);
        y_4 : out STD_LOGIC_VECTOR(15 downto 0);
        y_5 : out STD_LOGIC_VECTOR(15 downto 0);
        y_6 : out STD_LOGIC_VECTOR(15 downto 0);
        y_7 : out STD_LOGIC_VECTOR(15 downto 0);
        y_8 : out STD_LOGIC_VECTOR(15 downto 0);
        y_9 : out STD_LOGIC_VECTOR(15 downto 0);
        y_10 : out STD_LOGIC_VECTOR(15 downto 0);
        y_11 : out STD_LOGIC_VECTOR(15 downto 0);
        y_12 : out STD_LOGIC_VECTOR(15 downto 0);
        y_13 : out STD_LOGIC_VECTOR(15 downto 0);
        y_14 : out STD_LOGIC_VECTOR(15 downto 0);
        y_15 : out STD_LOGIC_VECTOR(15 downto 0);
        y_16 : out STD_LOGIC_VECTOR(15 downto 0);
        y_17 : out STD_LOGIC_VECTOR(15 downto 0);
        y_18 : out STD_LOGIC_VECTOR(15 downto 0);
        y_19 : out STD_LOGIC_VECTOR(15 downto 0);
        y_20 : out STD_LOGIC_VECTOR(15 downto 0);
        y_21 : out STD_LOGIC_VECTOR(15 downto 0);
        y_22 : out STD_LOGIC_VECTOR(15 downto 0);
        y_23 : out STD_LOGIC_VECTOR(15 downto 0);
        y_24 : out STD_LOGIC_VECTOR(15 downto 0);
        y_25 : out STD_LOGIC_VECTOR(15 downto 0);
        y_26 : out STD_LOGIC_VECTOR(15 downto 0);
        y_27 : out STD_LOGIC_VECTOR(15 downto 0);
        y_28 : out STD_LOGIC_VECTOR(15 downto 0);
        y_29 : out STD_LOGIC_VECTOR(15 downto 0);
        y_30 : out STD_LOGIC_VECTOR(15 downto 0);
        y_31 : out STD_LOGIC_VECTOR(15 downto 0);
        y_32 : out STD_LOGIC_VECTOR(15 downto 0);
        y_33 : out STD_LOGIC_VECTOR(15 downto 0);
        y_34 : out STD_LOGIC_VECTOR(15 downto 0);
        y_35 : out STD_LOGIC_VECTOR(15 downto 0);
        y_36 : out STD_LOGIC_VECTOR(15 downto 0);
        y_37 : out STD_LOGIC_VECTOR(15 downto 0);
        y_38 : out STD_LOGIC_VECTOR(15 downto 0);
        y_39 : out STD_LOGIC_VECTOR(15 downto 0);
        y_40 : out STD_LOGIC_VECTOR(15 downto 0);
        y_41 : out STD_LOGIC_VECTOR(15 downto 0);
        y_42 : out STD_LOGIC_VECTOR(15 downto 0);
        y_43 : out STD_LOGIC_VECTOR(15 downto 0);
        y_44 : out STD_LOGIC_VECTOR(15 downto 0);
        y_45 : out STD_LOGIC_VECTOR(15 downto 0);
        y_46 : out STD_LOGIC_VECTOR(15 downto 0);
        y_47 : out STD_LOGIC_VECTOR(15 downto 0);
        y_48 : out STD_LOGIC_VECTOR(15 downto 0);
        y_49 : out STD_LOGIC_VECTOR(15 downto 0);
        y_50 : out STD_LOGIC_VECTOR(15 downto 0);
        y_51 : out STD_LOGIC_VECTOR(15 downto 0);
        y_52 : out STD_LOGIC_VECTOR(15 downto 0);
        y_53 : out STD_LOGIC_VECTOR(15 downto 0);
        y_54 : out STD_LOGIC_VECTOR(15 downto 0);
        y_55 : out STD_LOGIC_VECTOR(15 downto 0);
        y_56 : out STD_LOGIC_VECTOR(15 downto 0);
        y_57 : out STD_LOGIC_VECTOR(15 downto 0);
        y_58 : out STD_LOGIC_VECTOR(15 downto 0);
        y_59 : out STD_LOGIC_VECTOR(15 downto 0);
        y_60 : out STD_LOGIC_VECTOR(15 downto 0);
        y_61 : out STD_LOGIC_VECTOR(15 downto 0);
        y_62 : out STD_LOGIC_VECTOR(15 downto 0);
        y_63 : out STD_LOGIC_VECTOR(15 downto 0);
        y_64 : out STD_LOGIC_VECTOR(15 downto 0);
        y_65 : out STD_LOGIC_VECTOR(15 downto 0);
        y_66 : out STD_LOGIC_VECTOR(15 downto 0);
        y_67 : out STD_LOGIC_VECTOR(15 downto 0);
        y_68 : out STD_LOGIC_VECTOR(15 downto 0);
        y_69 : out STD_LOGIC_VECTOR(15 downto 0);
        y_70 : out STD_LOGIC_VECTOR(15 downto 0);
        y_71 : out STD_LOGIC_VECTOR(15 downto 0);
        y_72 : out STD_LOGIC_VECTOR(15 downto 0);
        y_73 : out STD_LOGIC_VECTOR(15 downto 0);
        y_74 : out STD_LOGIC_VECTOR(15 downto 0);
        y_75 : out STD_LOGIC_VECTOR(15 downto 0);
        y_76 : out STD_LOGIC_VECTOR(15 downto 0);
        y_77 : out STD_LOGIC_VECTOR(15 downto 0);
        y_78 : out STD_LOGIC_VECTOR(15 downto 0);
        y_79 : out STD_LOGIC_VECTOR(15 downto 0);
        y_80 : out STD_LOGIC_VECTOR(15 downto 0);
        y_81 : out STD_LOGIC_VECTOR(15 downto 0);
        y_82 : out STD_LOGIC_VECTOR(15 downto 0);
        y_83 : out STD_LOGIC_VECTOR(15 downto 0);
        y_84 : out STD_LOGIC_VECTOR(15 downto 0);
        y_85 : out STD_LOGIC_VECTOR(15 downto 0);
        y_86 : out STD_LOGIC_VECTOR(15 downto 0);
        y_87 : out STD_LOGIC_VECTOR(15 downto 0);
        y_88 : out STD_LOGIC_VECTOR(15 downto 0);
        y_89 : out STD_LOGIC_VECTOR(15 downto 0);
        y_90 : out STD_LOGIC_VECTOR(15 downto 0);
        y_91 : out STD_LOGIC_VECTOR(15 downto 0);
        y_92 : out STD_LOGIC_VECTOR(15 downto 0);
        y_93 : out STD_LOGIC_VECTOR(15 downto 0);
        y_94 : out STD_LOGIC_VECTOR(15 downto 0);
        y_95 : out STD_LOGIC_VECTOR(15 downto 0);
        y_96 : out STD_LOGIC_VECTOR(15 downto 0);
        y_97 : out STD_LOGIC_VECTOR(15 downto 0);
        y_98 : out STD_LOGIC_VECTOR(15 downto 0);
        y_99 : out STD_LOGIC_VECTOR(15 downto 0);
        y_100 : out STD_LOGIC_VECTOR(15 downto 0);
        y_101 : out STD_LOGIC_VECTOR(15 downto 0);
        y_102 : out STD_LOGIC_VECTOR(15 downto 0);
        y_103 : out STD_LOGIC_VECTOR(15 downto 0);
        y_104 : out STD_LOGIC_VECTOR(15 downto 0);
        y_105 : out STD_LOGIC_VECTOR(15 downto 0);
        y_106 : out STD_LOGIC_VECTOR(15 downto 0);
        y_107 : out STD_LOGIC_VECTOR(15 downto 0);
        y_108 : out STD_LOGIC_VECTOR(15 downto 0);
        y_109 : out STD_LOGIC_VECTOR(15 downto 0);
        y_110 : out STD_LOGIC_VECTOR(15 downto 0);
        y_111 : out STD_LOGIC_VECTOR(15 downto 0);
        y_112 : out STD_LOGIC_VECTOR(15 downto 0);
        y_113 : out STD_LOGIC_VECTOR(15 downto 0);
        y_114 : out STD_LOGIC_VECTOR(15 downto 0);
        y_115 : out STD_LOGIC_VECTOR(15 downto 0);
        y_116 : out STD_LOGIC_VECTOR(15 downto 0);
        y_117 : out STD_LOGIC_VECTOR(15 downto 0);
        y_118 : out STD_LOGIC_VECTOR(15 downto 0);
        y_119 : out STD_LOGIC_VECTOR(15 downto 0);
        y_120 : out STD_LOGIC_VECTOR(15 downto 0);
        y_121 : out STD_LOGIC_VECTOR(15 downto 0);
        y_122 : out STD_LOGIC_VECTOR(15 downto 0);
        y_123 : out STD_LOGIC_VECTOR(15 downto 0);
        y_124 : out STD_LOGIC_VECTOR(15 downto 0);
        y_125 : out STD_LOGIC_VECTOR(15 downto 0);
        y_126 : out STD_LOGIC_VECTOR(15 downto 0);
        y_127 : out STD_LOGIC_VECTOR(15 downto 0);
        y_128 : out STD_LOGIC_VECTOR(15 downto 0);
        y_129 : out STD_LOGIC_VECTOR(15 downto 0);
        y_130 : out STD_LOGIC_VECTOR(15 downto 0);
        y_131 : out STD_LOGIC_VECTOR(15 downto 0);
        y_132 : out STD_LOGIC_VECTOR(15 downto 0);
        y_133 : out STD_LOGIC_VECTOR(15 downto 0);
        y_134 : out STD_LOGIC_VECTOR(15 downto 0);
        y_135 : out STD_LOGIC_VECTOR(15 downto 0);
        y_136 : out STD_LOGIC_VECTOR(15 downto 0);
        y_137 : out STD_LOGIC_VECTOR(15 downto 0);
        y_138 : out STD_LOGIC_VECTOR(15 downto 0);
        y_139 : out STD_LOGIC_VECTOR(15 downto 0);
        y_140 : out STD_LOGIC_VECTOR(15 downto 0);
        y_141 : out STD_LOGIC_VECTOR(15 downto 0);
        y_142 : out STD_LOGIC_VECTOR(15 downto 0);
        y_143 : out STD_LOGIC_VECTOR(15 downto 0);
        y_144 : out STD_LOGIC_VECTOR(15 downto 0);
        y_145 : out STD_LOGIC_VECTOR(15 downto 0);
        y_146 : out STD_LOGIC_VECTOR(15 downto 0);
        y_147 : out STD_LOGIC_VECTOR(15 downto 0);
        y_148 : out STD_LOGIC_VECTOR(15 downto 0);
        y_149 : out STD_LOGIC_VECTOR(15 downto 0);
        y_150 : out STD_LOGIC_VECTOR(15 downto 0);
        y_151 : out STD_LOGIC_VECTOR(15 downto 0);
        y_152 : out STD_LOGIC_VECTOR(15 downto 0);
        y_153 : out STD_LOGIC_VECTOR(15 downto 0);
        y_154 : out STD_LOGIC_VECTOR(15 downto 0);
        y_155 : out STD_LOGIC_VECTOR(15 downto 0);
        y_156 : out STD_LOGIC_VECTOR(15 downto 0);
        y_157 : out STD_LOGIC_VECTOR(15 downto 0);
        y_158 : out STD_LOGIC_VECTOR(15 downto 0);
        y_159 : out STD_LOGIC_VECTOR(15 downto 0);
        y_160 : out STD_LOGIC_VECTOR(15 downto 0);
        y_161 : out STD_LOGIC_VECTOR(15 downto 0);
        y_162 : out STD_LOGIC_VECTOR(15 downto 0);
        y_163 : out STD_LOGIC_VECTOR(15 downto 0);
        y_164 : out STD_LOGIC_VECTOR(15 downto 0);
        y_165 : out STD_LOGIC_VECTOR(15 downto 0);
        y_166 : out STD_LOGIC_VECTOR(15 downto 0);
        y_167 : out STD_LOGIC_VECTOR(15 downto 0);
        y_168 : out STD_LOGIC_VECTOR(15 downto 0);
        y_169 : out STD_LOGIC_VECTOR(15 downto 0);
        y_170 : out STD_LOGIC_VECTOR(15 downto 0);
        y_171 : out STD_LOGIC_VECTOR(15 downto 0);
        y_172 : out STD_LOGIC_VECTOR(15 downto 0);
        y_173 : out STD_LOGIC_VECTOR(15 downto 0);
        y_174 : out STD_LOGIC_VECTOR(15 downto 0);
        y_175 : out STD_LOGIC_VECTOR(15 downto 0);
        y_176 : out STD_LOGIC_VECTOR(15 downto 0);
        y_177 : out STD_LOGIC_VECTOR(15 downto 0);
        y_178 : out STD_LOGIC_VECTOR(15 downto 0);
        y_179 : out STD_LOGIC_VECTOR(15 downto 0);
        y_180 : out STD_LOGIC_VECTOR(15 downto 0);
        y_181 : out STD_LOGIC_VECTOR(15 downto 0);
        y_182 : out STD_LOGIC_VECTOR(15 downto 0);
        y_183 : out STD_LOGIC_VECTOR(15 downto 0);
        y_184 : out STD_LOGIC_VECTOR(15 downto 0);
        y_185 : out STD_LOGIC_VECTOR(15 downto 0);
        y_186 : out STD_LOGIC_VECTOR(15 downto 0);
        y_187 : out STD_LOGIC_VECTOR(15 downto 0);
        y_188 : out STD_LOGIC_VECTOR(15 downto 0);
        y_189 : out STD_LOGIC_VECTOR(15 downto 0);
        y_190 : out STD_LOGIC_VECTOR(15 downto 0);
        y_191 : out STD_LOGIC_VECTOR(15 downto 0);
        y_192 : out STD_LOGIC_VECTOR(15 downto 0);
        y_193 : out STD_LOGIC_VECTOR(15 downto 0);
        y_194 : out STD_LOGIC_VECTOR(15 downto 0);
        y_195 : out STD_LOGIC_VECTOR(15 downto 0);
        y_196 : out STD_LOGIC_VECTOR(15 downto 0);
        y_197 : out STD_LOGIC_VECTOR(15 downto 0);
        y_198 : out STD_LOGIC_VECTOR(15 downto 0);
        y_199 : out STD_LOGIC_VECTOR(15 downto 0);
        y_200 : out STD_LOGIC_VECTOR(15 downto 0);
        y_201 : out STD_LOGIC_VECTOR(15 downto 0);
        y_202 : out STD_LOGIC_VECTOR(15 downto 0);
        y_203 : out STD_LOGIC_VECTOR(15 downto 0);
        y_204 : out STD_LOGIC_VECTOR(15 downto 0);
        y_205 : out STD_LOGIC_VECTOR(15 downto 0);
        y_206 : out STD_LOGIC_VECTOR(15 downto 0);
        y_207 : out STD_LOGIC_VECTOR(15 downto 0);
        y_208 : out STD_LOGIC_VECTOR(15 downto 0);
        y_209 : out STD_LOGIC_VECTOR(15 downto 0);
        y_210 : out STD_LOGIC_VECTOR(15 downto 0);
        y_211 : out STD_LOGIC_VECTOR(15 downto 0);
        y_212 : out STD_LOGIC_VECTOR(15 downto 0);
        y_213 : out STD_LOGIC_VECTOR(15 downto 0);
        y_214 : out STD_LOGIC_VECTOR(15 downto 0);
        y_215 : out STD_LOGIC_VECTOR(15 downto 0);
        y_216 : out STD_LOGIC_VECTOR(15 downto 0);
        y_217 : out STD_LOGIC_VECTOR(15 downto 0);
        y_218 : out STD_LOGIC_VECTOR(15 downto 0);
        y_219 : out STD_LOGIC_VECTOR(15 downto 0);
        y_220 : out STD_LOGIC_VECTOR(15 downto 0);
        y_221 : out STD_LOGIC_VECTOR(15 downto 0);
        y_222 : out STD_LOGIC_VECTOR(15 downto 0);
        y_223 : out STD_LOGIC_VECTOR(15 downto 0);
        y_224 : out STD_LOGIC_VECTOR(15 downto 0);
        y_225 : out STD_LOGIC_VECTOR(15 downto 0);
        y_226 : out STD_LOGIC_VECTOR(15 downto 0);
        y_227 : out STD_LOGIC_VECTOR(15 downto 0);
        y_228 : out STD_LOGIC_VECTOR(15 downto 0);
        y_229 : out STD_LOGIC_VECTOR(15 downto 0);
        y_230 : out STD_LOGIC_VECTOR(15 downto 0);
        y_231 : out STD_LOGIC_VECTOR(15 downto 0);
        y_232 : out STD_LOGIC_VECTOR(15 downto 0);
        y_233 : out STD_LOGIC_VECTOR(15 downto 0);
        y_234 : out STD_LOGIC_VECTOR(15 downto 0);
        y_235 : out STD_LOGIC_VECTOR(15 downto 0);
        y_236 : out STD_LOGIC_VECTOR(15 downto 0);
        y_237 : out STD_LOGIC_VECTOR(15 downto 0);
        y_238 : out STD_LOGIC_VECTOR(15 downto 0);
        y_239 : out STD_LOGIC_VECTOR(15 downto 0);
        y_240 : out STD_LOGIC_VECTOR(15 downto 0);
        y_241 : out STD_LOGIC_VECTOR(15 downto 0);
        y_242 : out STD_LOGIC_VECTOR(15 downto 0);
        y_243 : out STD_LOGIC_VECTOR(15 downto 0);
        y_244 : out STD_LOGIC_VECTOR(15 downto 0);
        y_245 : out STD_LOGIC_VECTOR(15 downto 0);
        y_246 : out STD_LOGIC_VECTOR(15 downto 0);
        y_247 : out STD_LOGIC_VECTOR(15 downto 0);
        y_248 : out STD_LOGIC_VECTOR(15 downto 0);
        y_249 : out STD_LOGIC_VECTOR(15 downto 0);
        y_250 : out STD_LOGIC_VECTOR(15 downto 0);
        y_251 : out STD_LOGIC_VECTOR(15 downto 0);
        y_252 : out STD_LOGIC_VECTOR(15 downto 0);
        y_253 : out STD_LOGIC_VECTOR(15 downto 0);
        y_254 : out STD_LOGIC_VECTOR(15 downto 0);
        y_255 : out STD_LOGIC_VECTOR(15 downto 0);
        y_256 : out STD_LOGIC_VECTOR(15 downto 0);
        y_257 : out STD_LOGIC_VECTOR(15 downto 0);
        y_258 : out STD_LOGIC_VECTOR(15 downto 0);
        y_259 : out STD_LOGIC_VECTOR(15 downto 0);
        y_260 : out STD_LOGIC_VECTOR(15 downto 0);
        y_261 : out STD_LOGIC_VECTOR(15 downto 0);
        y_262 : out STD_LOGIC_VECTOR(15 downto 0);
        y_263 : out STD_LOGIC_VECTOR(15 downto 0);
        y_264 : out STD_LOGIC_VECTOR(15 downto 0);
        y_265 : out STD_LOGIC_VECTOR(15 downto 0);
        y_266 : out STD_LOGIC_VECTOR(15 downto 0);
        y_267 : out STD_LOGIC_VECTOR(15 downto 0);
        y_268 : out STD_LOGIC_VECTOR(15 downto 0);
        y_269 : out STD_LOGIC_VECTOR(15 downto 0);
        y_270 : out STD_LOGIC_VECTOR(15 downto 0);
        y_271 : out STD_LOGIC_VECTOR(15 downto 0);
        y_272 : out STD_LOGIC_VECTOR(15 downto 0);
        y_273 : out STD_LOGIC_VECTOR(15 downto 0);
        y_274 : out STD_LOGIC_VECTOR(15 downto 0);
        y_275 : out STD_LOGIC_VECTOR(15 downto 0);
        y_276 : out STD_LOGIC_VECTOR(15 downto 0);
        y_277 : out STD_LOGIC_VECTOR(15 downto 0);
        y_278 : out STD_LOGIC_VECTOR(15 downto 0);
        y_279 : out STD_LOGIC_VECTOR(15 downto 0);
        y_280 : out STD_LOGIC_VECTOR(15 downto 0);
        y_281 : out STD_LOGIC_VECTOR(15 downto 0);
        y_282 : out STD_LOGIC_VECTOR(15 downto 0);
        y_283 : out STD_LOGIC_VECTOR(15 downto 0);
        y_284 : out STD_LOGIC_VECTOR(15 downto 0);
        y_285 : out STD_LOGIC_VECTOR(15 downto 0);
        y_286 : out STD_LOGIC_VECTOR(15 downto 0);
        y_287 : out STD_LOGIC_VECTOR(15 downto 0);
        y_288 : out STD_LOGIC_VECTOR(15 downto 0);
        y_289 : out STD_LOGIC_VECTOR(15 downto 0);
        y_290 : out STD_LOGIC_VECTOR(15 downto 0);
        y_291 : out STD_LOGIC_VECTOR(15 downto 0);
        y_292 : out STD_LOGIC_VECTOR(15 downto 0);
        y_293 : out STD_LOGIC_VECTOR(15 downto 0);
        y_294 : out STD_LOGIC_VECTOR(15 downto 0);
        y_295 : out STD_LOGIC_VECTOR(15 downto 0);
        y_296 : out STD_LOGIC_VECTOR(15 downto 0);
        y_297 : out STD_LOGIC_VECTOR(15 downto 0);
        y_298 : out STD_LOGIC_VECTOR(15 downto 0);
        y_299 : out STD_LOGIC_VECTOR(15 downto 0);
        y_300 : out STD_LOGIC_VECTOR(15 downto 0);
        y_301 : out STD_LOGIC_VECTOR(15 downto 0);
        y_302 : out STD_LOGIC_VECTOR(15 downto 0);
        y_303 : out STD_LOGIC_VECTOR(15 downto 0);
        y_304 : out STD_LOGIC_VECTOR(15 downto 0);
        y_305 : out STD_LOGIC_VECTOR(15 downto 0);
        y_306 : out STD_LOGIC_VECTOR(15 downto 0);
        y_307 : out STD_LOGIC_VECTOR(15 downto 0);
        y_308 : out STD_LOGIC_VECTOR(15 downto 0);
        y_309 : out STD_LOGIC_VECTOR(15 downto 0);
        y_310 : out STD_LOGIC_VECTOR(15 downto 0);
        y_311 : out STD_LOGIC_VECTOR(15 downto 0);
        y_312 : out STD_LOGIC_VECTOR(15 downto 0);
        y_313 : out STD_LOGIC_VECTOR(15 downto 0);
        y_314 : out STD_LOGIC_VECTOR(15 downto 0);
        y_315 : out STD_LOGIC_VECTOR(15 downto 0);
        y_316 : out STD_LOGIC_VECTOR(15 downto 0);
        y_317 : out STD_LOGIC_VECTOR(15 downto 0);
        y_318 : out STD_LOGIC_VECTOR(15 downto 0);
        y_319 : out STD_LOGIC_VECTOR(15 downto 0);
        y_320 : out STD_LOGIC_VECTOR(15 downto 0);
        y_321 : out STD_LOGIC_VECTOR(15 downto 0);
        y_322 : out STD_LOGIC_VECTOR(15 downto 0);
        y_323 : out STD_LOGIC_VECTOR(15 downto 0);
        y_324 : out STD_LOGIC_VECTOR(15 downto 0);
        y_325 : out STD_LOGIC_VECTOR(15 downto 0);
        y_326 : out STD_LOGIC_VECTOR(15 downto 0);
        y_327 : out STD_LOGIC_VECTOR(15 downto 0);
        y_328 : out STD_LOGIC_VECTOR(15 downto 0);
        y_329 : out STD_LOGIC_VECTOR(15 downto 0);
        y_330 : out STD_LOGIC_VECTOR(15 downto 0);
        y_331 : out STD_LOGIC_VECTOR(15 downto 0);
        y_332 : out STD_LOGIC_VECTOR(15 downto 0);
        y_333 : out STD_LOGIC_VECTOR(15 downto 0);
        y_334 : out STD_LOGIC_VECTOR(15 downto 0);
        y_335 : out STD_LOGIC_VECTOR(15 downto 0);
        y_336 : out STD_LOGIC_VECTOR(15 downto 0);
        y_337 : out STD_LOGIC_VECTOR(15 downto 0);
        y_338 : out STD_LOGIC_VECTOR(15 downto 0);
        y_339 : out STD_LOGIC_VECTOR(15 downto 0);
        y_340 : out STD_LOGIC_VECTOR(15 downto 0);
        y_341 : out STD_LOGIC_VECTOR(15 downto 0);
        y_342 : out STD_LOGIC_VECTOR(15 downto 0);
        y_343 : out STD_LOGIC_VECTOR(15 downto 0);
        y_344 : out STD_LOGIC_VECTOR(15 downto 0);
        y_345 : out STD_LOGIC_VECTOR(15 downto 0);
        y_346 : out STD_LOGIC_VECTOR(15 downto 0);
        y_347 : out STD_LOGIC_VECTOR(15 downto 0);
        y_348 : out STD_LOGIC_VECTOR(15 downto 0);
        y_349 : out STD_LOGIC_VECTOR(15 downto 0);
        y_350 : out STD_LOGIC_VECTOR(15 downto 0);
        y_351 : out STD_LOGIC_VECTOR(15 downto 0);
        y_352 : out STD_LOGIC_VECTOR(15 downto 0);
        y_353 : out STD_LOGIC_VECTOR(15 downto 0);
        y_354 : out STD_LOGIC_VECTOR(15 downto 0);
        y_355 : out STD_LOGIC_VECTOR(15 downto 0);
        y_356 : out STD_LOGIC_VECTOR(15 downto 0);
        y_357 : out STD_LOGIC_VECTOR(15 downto 0);
        y_358 : out STD_LOGIC_VECTOR(15 downto 0);
        y_359 : out STD_LOGIC_VECTOR(15 downto 0);
        y_360 : out STD_LOGIC_VECTOR(15 downto 0);
        y_361 : out STD_LOGIC_VECTOR(15 downto 0);
        y_362 : out STD_LOGIC_VECTOR(15 downto 0);
        y_363 : out STD_LOGIC_VECTOR(15 downto 0);
        y_364 : out STD_LOGIC_VECTOR(15 downto 0);
        y_365 : out STD_LOGIC_VECTOR(15 downto 0);
        y_366 : out STD_LOGIC_VECTOR(15 downto 0);
        y_367 : out STD_LOGIC_VECTOR(15 downto 0);
        y_368 : out STD_LOGIC_VECTOR(15 downto 0);
        y_369 : out STD_LOGIC_VECTOR(15 downto 0);
        y_370 : out STD_LOGIC_VECTOR(15 downto 0);
        y_371 : out STD_LOGIC_VECTOR(15 downto 0);
        y_372 : out STD_LOGIC_VECTOR(15 downto 0);
        y_373 : out STD_LOGIC_VECTOR(15 downto 0);
        y_374 : out STD_LOGIC_VECTOR(15 downto 0);
        y_375 : out STD_LOGIC_VECTOR(15 downto 0);
        y_376 : out STD_LOGIC_VECTOR(15 downto 0);
        y_377 : out STD_LOGIC_VECTOR(15 downto 0);
        y_378 : out STD_LOGIC_VECTOR(15 downto 0);
        y_379 : out STD_LOGIC_VECTOR(15 downto 0);
        y_380 : out STD_LOGIC_VECTOR(15 downto 0);
        y_381 : out STD_LOGIC_VECTOR(15 downto 0);
        y_382 : out STD_LOGIC_VECTOR(15 downto 0);
        y_383 : out STD_LOGIC_VECTOR(15 downto 0);
        y_384 : out STD_LOGIC_VECTOR(15 downto 0);
        y_385 : out STD_LOGIC_VECTOR(15 downto 0);
        y_386 : out STD_LOGIC_VECTOR(15 downto 0);
        y_387 : out STD_LOGIC_VECTOR(15 downto 0);
        y_388 : out STD_LOGIC_VECTOR(15 downto 0);
        y_389 : out STD_LOGIC_VECTOR(15 downto 0);
        y_390 : out STD_LOGIC_VECTOR(15 downto 0);
        y_391 : out STD_LOGIC_VECTOR(15 downto 0);
        y_392 : out STD_LOGIC_VECTOR(15 downto 0);
        y_393 : out STD_LOGIC_VECTOR(15 downto 0);
        y_394 : out STD_LOGIC_VECTOR(15 downto 0);
        y_395 : out STD_LOGIC_VECTOR(15 downto 0);
        y_396 : out STD_LOGIC_VECTOR(15 downto 0);
        y_397 : out STD_LOGIC_VECTOR(15 downto 0);
        y_398 : out STD_LOGIC_VECTOR(15 downto 0);
        y_399 : out STD_LOGIC_VECTOR(15 downto 0);
        y_400 : out STD_LOGIC_VECTOR(15 downto 0);
        y_401 : out STD_LOGIC_VECTOR(15 downto 0);
        y_402 : out STD_LOGIC_VECTOR(15 downto 0);
        y_403 : out STD_LOGIC_VECTOR(15 downto 0);
        y_404 : out STD_LOGIC_VECTOR(15 downto 0);
        y_405 : out STD_LOGIC_VECTOR(15 downto 0);
        y_406 : out STD_LOGIC_VECTOR(15 downto 0);
        y_407 : out STD_LOGIC_VECTOR(15 downto 0);
        y_408 : out STD_LOGIC_VECTOR(15 downto 0);
        y_409 : out STD_LOGIC_VECTOR(15 downto 0);
        y_410 : out STD_LOGIC_VECTOR(15 downto 0);
        y_411 : out STD_LOGIC_VECTOR(15 downto 0);
        y_412 : out STD_LOGIC_VECTOR(15 downto 0);
        y_413 : out STD_LOGIC_VECTOR(15 downto 0);
        y_414 : out STD_LOGIC_VECTOR(15 downto 0);
        y_415 : out STD_LOGIC_VECTOR(15 downto 0);
        y_416 : out STD_LOGIC_VECTOR(15 downto 0);
        y_417 : out STD_LOGIC_VECTOR(15 downto 0);
        y_418 : out STD_LOGIC_VECTOR(15 downto 0);
        y_419 : out STD_LOGIC_VECTOR(15 downto 0);
        y_420 : out STD_LOGIC_VECTOR(15 downto 0);
        y_421 : out STD_LOGIC_VECTOR(15 downto 0);
        y_422 : out STD_LOGIC_VECTOR(15 downto 0);
        y_423 : out STD_LOGIC_VECTOR(15 downto 0);
        y_424 : out STD_LOGIC_VECTOR(15 downto 0);
        y_425 : out STD_LOGIC_VECTOR(15 downto 0);
        y_426 : out STD_LOGIC_VECTOR(15 downto 0);
        y_427 : out STD_LOGIC_VECTOR(15 downto 0);
        y_428 : out STD_LOGIC_VECTOR(15 downto 0);
        y_429 : out STD_LOGIC_VECTOR(15 downto 0);
        y_430 : out STD_LOGIC_VECTOR(15 downto 0);
        y_431 : out STD_LOGIC_VECTOR(15 downto 0);
        y_432 : out STD_LOGIC_VECTOR(15 downto 0);
        y_433 : out STD_LOGIC_VECTOR(15 downto 0);
        y_434 : out STD_LOGIC_VECTOR(15 downto 0);
        y_435 : out STD_LOGIC_VECTOR(15 downto 0);
        y_436 : out STD_LOGIC_VECTOR(15 downto 0);
        y_437 : out STD_LOGIC_VECTOR(15 downto 0);
        y_438 : out STD_LOGIC_VECTOR(15 downto 0);
        y_439 : out STD_LOGIC_VECTOR(15 downto 0);
        y_440 : out STD_LOGIC_VECTOR(15 downto 0);
        y_441 : out STD_LOGIC_VECTOR(15 downto 0);
        y_442 : out STD_LOGIC_VECTOR(15 downto 0);
        y_443 : out STD_LOGIC_VECTOR(15 downto 0);
        y_444 : out STD_LOGIC_VECTOR(15 downto 0);
        y_445 : out STD_LOGIC_VECTOR(15 downto 0);
        y_446 : out STD_LOGIC_VECTOR(15 downto 0);
        y_447 : out STD_LOGIC_VECTOR(15 downto 0);
        y_448 : out STD_LOGIC_VECTOR(15 downto 0);
        y_449 : out STD_LOGIC_VECTOR(15 downto 0);
        y_450 : out STD_LOGIC_VECTOR(15 downto 0);
        y_451 : out STD_LOGIC_VECTOR(15 downto 0);
        y_452 : out STD_LOGIC_VECTOR(15 downto 0);
        y_453 : out STD_LOGIC_VECTOR(15 downto 0);
        y_454 : out STD_LOGIC_VECTOR(15 downto 0);
        y_455 : out STD_LOGIC_VECTOR(15 downto 0);
        y_456 : out STD_LOGIC_VECTOR(15 downto 0);
        y_457 : out STD_LOGIC_VECTOR(15 downto 0);
        y_458 : out STD_LOGIC_VECTOR(15 downto 0);
        y_459 : out STD_LOGIC_VECTOR(15 downto 0);
        y_460 : out STD_LOGIC_VECTOR(15 downto 0);
        y_461 : out STD_LOGIC_VECTOR(15 downto 0);
        y_462 : out STD_LOGIC_VECTOR(15 downto 0);
        y_463 : out STD_LOGIC_VECTOR(15 downto 0);
        y_464 : out STD_LOGIC_VECTOR(15 downto 0);
        y_465 : out STD_LOGIC_VECTOR(15 downto 0);
        y_466 : out STD_LOGIC_VECTOR(15 downto 0);
        y_467 : out STD_LOGIC_VECTOR(15 downto 0);
        y_468 : out STD_LOGIC_VECTOR(15 downto 0);
        y_469 : out STD_LOGIC_VECTOR(15 downto 0);
        y_470 : out STD_LOGIC_VECTOR(15 downto 0);
        y_471 : out STD_LOGIC_VECTOR(15 downto 0);
        y_472 : out STD_LOGIC_VECTOR(15 downto 0);
        y_473 : out STD_LOGIC_VECTOR(15 downto 0);
        y_474 : out STD_LOGIC_VECTOR(15 downto 0);
        y_475 : out STD_LOGIC_VECTOR(15 downto 0);
        y_476 : out STD_LOGIC_VECTOR(15 downto 0);
        y_477 : out STD_LOGIC_VECTOR(15 downto 0);
        y_478 : out STD_LOGIC_VECTOR(15 downto 0);
        y_479 : out STD_LOGIC_VECTOR(15 downto 0);
        y_480 : out STD_LOGIC_VECTOR(15 downto 0);
        y_481 : out STD_LOGIC_VECTOR(15 downto 0);
        y_482 : out STD_LOGIC_VECTOR(15 downto 0);
        y_483 : out STD_LOGIC_VECTOR(15 downto 0);
        y_484 : out STD_LOGIC_VECTOR(15 downto 0);
        y_485 : out STD_LOGIC_VECTOR(15 downto 0);
        y_486 : out STD_LOGIC_VECTOR(15 downto 0);
        y_487 : out STD_LOGIC_VECTOR(15 downto 0);
        y_488 : out STD_LOGIC_VECTOR(15 downto 0);
        y_489 : out STD_LOGIC_VECTOR(15 downto 0);
        y_490 : out STD_LOGIC_VECTOR(15 downto 0);
        y_491 : out STD_LOGIC_VECTOR(15 downto 0);
        y_492 : out STD_LOGIC_VECTOR(15 downto 0);
        y_493 : out STD_LOGIC_VECTOR(15 downto 0);
        y_494 : out STD_LOGIC_VECTOR(15 downto 0);
        y_495 : out STD_LOGIC_VECTOR(15 downto 0);
        y_496 : out STD_LOGIC_VECTOR(15 downto 0);
        y_497 : out STD_LOGIC_VECTOR(15 downto 0);
        y_498 : out STD_LOGIC_VECTOR(15 downto 0);
        y_499 : out STD_LOGIC_VECTOR(15 downto 0);
        y_500 : out STD_LOGIC_VECTOR(15 downto 0);
        y_501 : out STD_LOGIC_VECTOR(15 downto 0);
        y_502 : out STD_LOGIC_VECTOR(15 downto 0);
        y_503 : out STD_LOGIC_VECTOR(15 downto 0);
        y_504 : out STD_LOGIC_VECTOR(15 downto 0);
        y_505 : out STD_LOGIC_VECTOR(15 downto 0);
        y_506 : out STD_LOGIC_VECTOR(15 downto 0);
        y_507 : out STD_LOGIC_VECTOR(15 downto 0);
        y_508 : out STD_LOGIC_VECTOR(15 downto 0);
        y_509 : out STD_LOGIC_VECTOR(15 downto 0);
        y_510 : out STD_LOGIC_VECTOR(15 downto 0);
        y_511 : out STD_LOGIC_VECTOR(15 downto 0);
        y_512 : out STD_LOGIC_VECTOR(15 downto 0);
        y_513 : out STD_LOGIC_VECTOR(15 downto 0);
        y_514 : out STD_LOGIC_VECTOR(15 downto 0);
        y_515 : out STD_LOGIC_VECTOR(15 downto 0);
        y_516 : out STD_LOGIC_VECTOR(15 downto 0);
        y_517 : out STD_LOGIC_VECTOR(15 downto 0);
        y_518 : out STD_LOGIC_VECTOR(15 downto 0);
        y_519 : out STD_LOGIC_VECTOR(15 downto 0);
        y_520 : out STD_LOGIC_VECTOR(15 downto 0);
        y_521 : out STD_LOGIC_VECTOR(15 downto 0);
        y_522 : out STD_LOGIC_VECTOR(15 downto 0);
        y_523 : out STD_LOGIC_VECTOR(15 downto 0);
        y_524 : out STD_LOGIC_VECTOR(15 downto 0);
        y_525 : out STD_LOGIC_VECTOR(15 downto 0);
        y_526 : out STD_LOGIC_VECTOR(15 downto 0);
        y_527 : out STD_LOGIC_VECTOR(15 downto 0);
        y_528 : out STD_LOGIC_VECTOR(15 downto 0);
        y_529 : out STD_LOGIC_VECTOR(15 downto 0);
        y_530 : out STD_LOGIC_VECTOR(15 downto 0);
        y_531 : out STD_LOGIC_VECTOR(15 downto 0);
        y_532 : out STD_LOGIC_VECTOR(15 downto 0);
        y_533 : out STD_LOGIC_VECTOR(15 downto 0);
        y_534 : out STD_LOGIC_VECTOR(15 downto 0);
        y_535 : out STD_LOGIC_VECTOR(15 downto 0);
        y_536 : out STD_LOGIC_VECTOR(15 downto 0);
        y_537 : out STD_LOGIC_VECTOR(15 downto 0);
        y_538 : out STD_LOGIC_VECTOR(15 downto 0);
        y_539 : out STD_LOGIC_VECTOR(15 downto 0);
        y_540 : out STD_LOGIC_VECTOR(15 downto 0);
        y_541 : out STD_LOGIC_VECTOR(15 downto 0);
        y_542 : out STD_LOGIC_VECTOR(15 downto 0);
        y_543 : out STD_LOGIC_VECTOR(15 downto 0);
        y_544 : out STD_LOGIC_VECTOR(15 downto 0);
        y_545 : out STD_LOGIC_VECTOR(15 downto 0);
        y_546 : out STD_LOGIC_VECTOR(15 downto 0);
        y_547 : out STD_LOGIC_VECTOR(15 downto 0);
        y_548 : out STD_LOGIC_VECTOR(15 downto 0);
        y_549 : out STD_LOGIC_VECTOR(15 downto 0);
        y_550 : out STD_LOGIC_VECTOR(15 downto 0);
        y_551 : out STD_LOGIC_VECTOR(15 downto 0);
        y_552 : out STD_LOGIC_VECTOR(15 downto 0);
        y_553 : out STD_LOGIC_VECTOR(15 downto 0);
        y_554 : out STD_LOGIC_VECTOR(15 downto 0);
        y_555 : out STD_LOGIC_VECTOR(15 downto 0);
        y_556 : out STD_LOGIC_VECTOR(15 downto 0);
        y_557 : out STD_LOGIC_VECTOR(15 downto 0);
        y_558 : out STD_LOGIC_VECTOR(15 downto 0);
        y_559 : out STD_LOGIC_VECTOR(15 downto 0);
        y_560 : out STD_LOGIC_VECTOR(15 downto 0);
        y_561 : out STD_LOGIC_VECTOR(15 downto 0);
        y_562 : out STD_LOGIC_VECTOR(15 downto 0);
        y_563 : out STD_LOGIC_VECTOR(15 downto 0);
        y_564 : out STD_LOGIC_VECTOR(15 downto 0);
        y_565 : out STD_LOGIC_VECTOR(15 downto 0);
        y_566 : out STD_LOGIC_VECTOR(15 downto 0);
        y_567 : out STD_LOGIC_VECTOR(15 downto 0);
        y_568 : out STD_LOGIC_VECTOR(15 downto 0);
        y_569 : out STD_LOGIC_VECTOR(15 downto 0);
        y_570 : out STD_LOGIC_VECTOR(15 downto 0);
        y_571 : out STD_LOGIC_VECTOR(15 downto 0);
        y_572 : out STD_LOGIC_VECTOR(15 downto 0);
        y_573 : out STD_LOGIC_VECTOR(15 downto 0);
        y_574 : out STD_LOGIC_VECTOR(15 downto 0);
        y_575 : out STD_LOGIC_VECTOR(15 downto 0);
        y_576 : out STD_LOGIC_VECTOR(15 downto 0);
        y_577 : out STD_LOGIC_VECTOR(15 downto 0);
        y_578 : out STD_LOGIC_VECTOR(15 downto 0);
        y_579 : out STD_LOGIC_VECTOR(15 downto 0);
        y_580 : out STD_LOGIC_VECTOR(15 downto 0);
        y_581 : out STD_LOGIC_VECTOR(15 downto 0);
        y_582 : out STD_LOGIC_VECTOR(15 downto 0);
        y_583 : out STD_LOGIC_VECTOR(15 downto 0);
        y_584 : out STD_LOGIC_VECTOR(15 downto 0);
        y_585 : out STD_LOGIC_VECTOR(15 downto 0);
        y_586 : out STD_LOGIC_VECTOR(15 downto 0);
        y_587 : out STD_LOGIC_VECTOR(15 downto 0);
        y_588 : out STD_LOGIC_VECTOR(15 downto 0);
        y_589 : out STD_LOGIC_VECTOR(15 downto 0);
        y_590 : out STD_LOGIC_VECTOR(15 downto 0);
        y_591 : out STD_LOGIC_VECTOR(15 downto 0);
        y_592 : out STD_LOGIC_VECTOR(15 downto 0);
        y_593 : out STD_LOGIC_VECTOR(15 downto 0);
        y_594 : out STD_LOGIC_VECTOR(15 downto 0);
        y_595 : out STD_LOGIC_VECTOR(15 downto 0);
        y_596 : out STD_LOGIC_VECTOR(15 downto 0);
        y_597 : out STD_LOGIC_VECTOR(15 downto 0);
        y_598 : out STD_LOGIC_VECTOR(15 downto 0);
        y_599 : out STD_LOGIC_VECTOR(15 downto 0);
        y_600 : out STD_LOGIC_VECTOR(15 downto 0);
        y_601 : out STD_LOGIC_VECTOR(15 downto 0);
        y_602 : out STD_LOGIC_VECTOR(15 downto 0);
        y_603 : out STD_LOGIC_VECTOR(15 downto 0);
        y_604 : out STD_LOGIC_VECTOR(15 downto 0);
        y_605 : out STD_LOGIC_VECTOR(15 downto 0);
        y_606 : out STD_LOGIC_VECTOR(15 downto 0);
        y_607 : out STD_LOGIC_VECTOR(15 downto 0);
        y_608 : out STD_LOGIC_VECTOR(15 downto 0);
        y_609 : out STD_LOGIC_VECTOR(15 downto 0);
        y_610 : out STD_LOGIC_VECTOR(15 downto 0);
        y_611 : out STD_LOGIC_VECTOR(15 downto 0);
        y_612 : out STD_LOGIC_VECTOR(15 downto 0);
        y_613 : out STD_LOGIC_VECTOR(15 downto 0);
        y_614 : out STD_LOGIC_VECTOR(15 downto 0);
        y_615 : out STD_LOGIC_VECTOR(15 downto 0);
        y_616 : out STD_LOGIC_VECTOR(15 downto 0);
        y_617 : out STD_LOGIC_VECTOR(15 downto 0);
        y_618 : out STD_LOGIC_VECTOR(15 downto 0);
        y_619 : out STD_LOGIC_VECTOR(15 downto 0);
        y_620 : out STD_LOGIC_VECTOR(15 downto 0);
        y_621 : out STD_LOGIC_VECTOR(15 downto 0);
        y_622 : out STD_LOGIC_VECTOR(15 downto 0);
        y_623 : out STD_LOGIC_VECTOR(15 downto 0);
        y_624 : out STD_LOGIC_VECTOR(15 downto 0);
        y_625 : out STD_LOGIC_VECTOR(15 downto 0);
        y_626 : out STD_LOGIC_VECTOR(15 downto 0);
        y_627 : out STD_LOGIC_VECTOR(15 downto 0);
        y_628 : out STD_LOGIC_VECTOR(15 downto 0);
        y_629 : out STD_LOGIC_VECTOR(15 downto 0);
        y_630 : out STD_LOGIC_VECTOR(15 downto 0);
        y_631 : out STD_LOGIC_VECTOR(15 downto 0);
        y_632 : out STD_LOGIC_VECTOR(15 downto 0);
        y_633 : out STD_LOGIC_VECTOR(15 downto 0);
        y_634 : out STD_LOGIC_VECTOR(15 downto 0);
        y_635 : out STD_LOGIC_VECTOR(15 downto 0);
        y_636 : out STD_LOGIC_VECTOR(15 downto 0);
        y_637 : out STD_LOGIC_VECTOR(15 downto 0);
        y_638 : out STD_LOGIC_VECTOR(15 downto 0);
        y_639 : out STD_LOGIC_VECTOR(15 downto 0);
        y_640 : out STD_LOGIC_VECTOR(15 downto 0);
        y_641 : out STD_LOGIC_VECTOR(15 downto 0);
        y_642 : out STD_LOGIC_VECTOR(15 downto 0);
        y_643 : out STD_LOGIC_VECTOR(15 downto 0);
        y_644 : out STD_LOGIC_VECTOR(15 downto 0);
        y_645 : out STD_LOGIC_VECTOR(15 downto 0);
        y_646 : out STD_LOGIC_VECTOR(15 downto 0);
        y_647 : out STD_LOGIC_VECTOR(15 downto 0);
        y_648 : out STD_LOGIC_VECTOR(15 downto 0);
        y_649 : out STD_LOGIC_VECTOR(15 downto 0);
        y_650 : out STD_LOGIC_VECTOR(15 downto 0);
        y_651 : out STD_LOGIC_VECTOR(15 downto 0);
        y_652 : out STD_LOGIC_VECTOR(15 downto 0);
        y_653 : out STD_LOGIC_VECTOR(15 downto 0);
        y_654 : out STD_LOGIC_VECTOR(15 downto 0);
        y_655 : out STD_LOGIC_VECTOR(15 downto 0);
        y_656 : out STD_LOGIC_VECTOR(15 downto 0);
        y_657 : out STD_LOGIC_VECTOR(15 downto 0);
        y_658 : out STD_LOGIC_VECTOR(15 downto 0);
        y_659 : out STD_LOGIC_VECTOR(15 downto 0);
        y_660 : out STD_LOGIC_VECTOR(15 downto 0);
        y_661 : out STD_LOGIC_VECTOR(15 downto 0);
        y_662 : out STD_LOGIC_VECTOR(15 downto 0);
        y_663 : out STD_LOGIC_VECTOR(15 downto 0);
        y_664 : out STD_LOGIC_VECTOR(15 downto 0);
        y_665 : out STD_LOGIC_VECTOR(15 downto 0);
        y_666 : out STD_LOGIC_VECTOR(15 downto 0);
        y_667 : out STD_LOGIC_VECTOR(15 downto 0);
        y_668 : out STD_LOGIC_VECTOR(15 downto 0);
        y_669 : out STD_LOGIC_VECTOR(15 downto 0);
        y_670 : out STD_LOGIC_VECTOR(15 downto 0);
        y_671 : out STD_LOGIC_VECTOR(15 downto 0);
        y_672 : out STD_LOGIC_VECTOR(15 downto 0);
        y_673 : out STD_LOGIC_VECTOR(15 downto 0);
        y_674 : out STD_LOGIC_VECTOR(15 downto 0);
        y_675 : out STD_LOGIC_VECTOR(15 downto 0);
        y_676 : out STD_LOGIC_VECTOR(15 downto 0);
        y_677 : out STD_LOGIC_VECTOR(15 downto 0);
        y_678 : out STD_LOGIC_VECTOR(15 downto 0);
        y_679 : out STD_LOGIC_VECTOR(15 downto 0);
        y_680 : out STD_LOGIC_VECTOR(15 downto 0);
        y_681 : out STD_LOGIC_VECTOR(15 downto 0);
        y_682 : out STD_LOGIC_VECTOR(15 downto 0);
        y_683 : out STD_LOGIC_VECTOR(15 downto 0);
        y_684 : out STD_LOGIC_VECTOR(15 downto 0);
        y_685 : out STD_LOGIC_VECTOR(15 downto 0);
        y_686 : out STD_LOGIC_VECTOR(15 downto 0);
        y_687 : out STD_LOGIC_VECTOR(15 downto 0);
        y_688 : out STD_LOGIC_VECTOR(15 downto 0);
        y_689 : out STD_LOGIC_VECTOR(15 downto 0);
        y_690 : out STD_LOGIC_VECTOR(15 downto 0);
        y_691 : out STD_LOGIC_VECTOR(15 downto 0);
        y_692 : out STD_LOGIC_VECTOR(15 downto 0);
        y_693 : out STD_LOGIC_VECTOR(15 downto 0);
        y_694 : out STD_LOGIC_VECTOR(15 downto 0);
        y_695 : out STD_LOGIC_VECTOR(15 downto 0);
        y_696 : out STD_LOGIC_VECTOR(15 downto 0);
        y_697 : out STD_LOGIC_VECTOR(15 downto 0);
        y_698 : out STD_LOGIC_VECTOR(15 downto 0);
        y_699 : out STD_LOGIC_VECTOR(15 downto 0);
        y_700 : out STD_LOGIC_VECTOR(15 downto 0);
        y_701 : out STD_LOGIC_VECTOR(15 downto 0);
        y_702 : out STD_LOGIC_VECTOR(15 downto 0);
        y_703 : out STD_LOGIC_VECTOR(15 downto 0);
        y_704 : out STD_LOGIC_VECTOR(15 downto 0);
        y_705 : out STD_LOGIC_VECTOR(15 downto 0);
        y_706 : out STD_LOGIC_VECTOR(15 downto 0);
        y_707 : out STD_LOGIC_VECTOR(15 downto 0);
        y_708 : out STD_LOGIC_VECTOR(15 downto 0);
        y_709 : out STD_LOGIC_VECTOR(15 downto 0);
        y_710 : out STD_LOGIC_VECTOR(15 downto 0);
        y_711 : out STD_LOGIC_VECTOR(15 downto 0);
        y_712 : out STD_LOGIC_VECTOR(15 downto 0);
        y_713 : out STD_LOGIC_VECTOR(15 downto 0);
        y_714 : out STD_LOGIC_VECTOR(15 downto 0);
        y_715 : out STD_LOGIC_VECTOR(15 downto 0);
        y_716 : out STD_LOGIC_VECTOR(15 downto 0);
        y_717 : out STD_LOGIC_VECTOR(15 downto 0);
        y_718 : out STD_LOGIC_VECTOR(15 downto 0);
        y_719 : out STD_LOGIC_VECTOR(15 downto 0);
        y_720 : out STD_LOGIC_VECTOR(15 downto 0);
        y_721 : out STD_LOGIC_VECTOR(15 downto 0);
        y_722 : out STD_LOGIC_VECTOR(15 downto 0);
        y_723 : out STD_LOGIC_VECTOR(15 downto 0);
        y_724 : out STD_LOGIC_VECTOR(15 downto 0);
        y_725 : out STD_LOGIC_VECTOR(15 downto 0);
        y_726 : out STD_LOGIC_VECTOR(15 downto 0);
        y_727 : out STD_LOGIC_VECTOR(15 downto 0);
        y_728 : out STD_LOGIC_VECTOR(15 downto 0);
        y_729 : out STD_LOGIC_VECTOR(15 downto 0);
        y_730 : out STD_LOGIC_VECTOR(15 downto 0);
        y_731 : out STD_LOGIC_VECTOR(15 downto 0);
        y_732 : out STD_LOGIC_VECTOR(15 downto 0);
        y_733 : out STD_LOGIC_VECTOR(15 downto 0);
        y_734 : out STD_LOGIC_VECTOR(15 downto 0);
        y_735 : out STD_LOGIC_VECTOR(15 downto 0);
        y_736 : out STD_LOGIC_VECTOR(15 downto 0);
        y_737 : out STD_LOGIC_VECTOR(15 downto 0);
        y_738 : out STD_LOGIC_VECTOR(15 downto 0);
        y_739 : out STD_LOGIC_VECTOR(15 downto 0);
        y_740 : out STD_LOGIC_VECTOR(15 downto 0);
        y_741 : out STD_LOGIC_VECTOR(15 downto 0);
        y_742 : out STD_LOGIC_VECTOR(15 downto 0);
        y_743 : out STD_LOGIC_VECTOR(15 downto 0);
        y_744 : out STD_LOGIC_VECTOR(15 downto 0);
        y_745 : out STD_LOGIC_VECTOR(15 downto 0);
        y_746 : out STD_LOGIC_VECTOR(15 downto 0);
        y_747 : out STD_LOGIC_VECTOR(15 downto 0);
        y_748 : out STD_LOGIC_VECTOR(15 downto 0);
        y_749 : out STD_LOGIC_VECTOR(15 downto 0);
        y_750 : out STD_LOGIC_VECTOR(15 downto 0);
        y_751 : out STD_LOGIC_VECTOR(15 downto 0);
        y_752 : out STD_LOGIC_VECTOR(15 downto 0);
        y_753 : out STD_LOGIC_VECTOR(15 downto 0);
        y_754 : out STD_LOGIC_VECTOR(15 downto 0);
        y_755 : out STD_LOGIC_VECTOR(15 downto 0);
        y_756 : out STD_LOGIC_VECTOR(15 downto 0);
        y_757 : out STD_LOGIC_VECTOR(15 downto 0);
        y_758 : out STD_LOGIC_VECTOR(15 downto 0);
        y_759 : out STD_LOGIC_VECTOR(15 downto 0);
        y_760 : out STD_LOGIC_VECTOR(15 downto 0);
        y_761 : out STD_LOGIC_VECTOR(15 downto 0);
        y_762 : out STD_LOGIC_VECTOR(15 downto 0);
        y_763 : out STD_LOGIC_VECTOR(15 downto 0);
        y_764 : out STD_LOGIC_VECTOR(15 downto 0);
        y_765 : out STD_LOGIC_VECTOR(15 downto 0);
        y_766 : out STD_LOGIC_VECTOR(15 downto 0);
        y_767 : out STD_LOGIC_VECTOR(15 downto 0);
        y_768 : out STD_LOGIC_VECTOR(15 downto 0);
        y_769 : out STD_LOGIC_VECTOR(15 downto 0);
        y_770 : out STD_LOGIC_VECTOR(15 downto 0);
        y_771 : out STD_LOGIC_VECTOR(15 downto 0);
        y_772 : out STD_LOGIC_VECTOR(15 downto 0);
        y_773 : out STD_LOGIC_VECTOR(15 downto 0);
        y_774 : out STD_LOGIC_VECTOR(15 downto 0);
        y_775 : out STD_LOGIC_VECTOR(15 downto 0);
        y_776 : out STD_LOGIC_VECTOR(15 downto 0);
        y_777 : out STD_LOGIC_VECTOR(15 downto 0);
        y_778 : out STD_LOGIC_VECTOR(15 downto 0);
        y_779 : out STD_LOGIC_VECTOR(15 downto 0);
        y_780 : out STD_LOGIC_VECTOR(15 downto 0);
        y_781 : out STD_LOGIC_VECTOR(15 downto 0);
        y_782 : out STD_LOGIC_VECTOR(15 downto 0);
	   y_783 : out STD_LOGIC_VECTOR(15 downto 0));
end component lstm_layer;

component  fully_connected_layer is
	Port (
		clk : in std_logic;
        x_0 : in STD_LOGIC_VECTOR(15 downto 0);
        x_1 : in STD_LOGIC_VECTOR(15 downto 0);
        x_2 : in STD_LOGIC_VECTOR(15 downto 0);
        x_3 : in STD_LOGIC_VECTOR(15 downto 0);
        x_4 : in STD_LOGIC_VECTOR(15 downto 0);
        x_5 : in STD_LOGIC_VECTOR(15 downto 0);
        x_6 : in STD_LOGIC_VECTOR(15 downto 0);
        x_7 : in STD_LOGIC_VECTOR(15 downto 0);
        x_8 : in STD_LOGIC_VECTOR(15 downto 0);
        x_9 : in STD_LOGIC_VECTOR(15 downto 0);
        x_10 : in STD_LOGIC_VECTOR(15 downto 0);
        x_11 : in STD_LOGIC_VECTOR(15 downto 0);
        x_12 : in STD_LOGIC_VECTOR(15 downto 0);
        x_13 : in STD_LOGIC_VECTOR(15 downto 0);
        x_14 : in STD_LOGIC_VECTOR(15 downto 0);
        x_15 : in STD_LOGIC_VECTOR(15 downto 0);
        x_16 : in STD_LOGIC_VECTOR(15 downto 0);
        x_17 : in STD_LOGIC_VECTOR(15 downto 0);
        x_18 : in STD_LOGIC_VECTOR(15 downto 0);
        x_19 : in STD_LOGIC_VECTOR(15 downto 0);
        x_20 : in STD_LOGIC_VECTOR(15 downto 0);
        x_21 : in STD_LOGIC_VECTOR(15 downto 0);
        x_22 : in STD_LOGIC_VECTOR(15 downto 0);
        x_23 : in STD_LOGIC_VECTOR(15 downto 0);
        x_24 : in STD_LOGIC_VECTOR(15 downto 0);
        x_25 : in STD_LOGIC_VECTOR(15 downto 0);
        x_26 : in STD_LOGIC_VECTOR(15 downto 0);
        x_27 : in STD_LOGIC_VECTOR(15 downto 0);
        x_28 : in STD_LOGIC_VECTOR(15 downto 0);
        x_29 : in STD_LOGIC_VECTOR(15 downto 0);
        x_30 : in STD_LOGIC_VECTOR(15 downto 0);
        x_31 : in STD_LOGIC_VECTOR(15 downto 0);
        x_32 : in STD_LOGIC_VECTOR(15 downto 0);
        x_33 : in STD_LOGIC_VECTOR(15 downto 0);
        x_34 : in STD_LOGIC_VECTOR(15 downto 0);
        x_35 : in STD_LOGIC_VECTOR(15 downto 0);
        x_36 : in STD_LOGIC_VECTOR(15 downto 0);
        x_37 : in STD_LOGIC_VECTOR(15 downto 0);
        x_38 : in STD_LOGIC_VECTOR(15 downto 0);
        x_39 : in STD_LOGIC_VECTOR(15 downto 0);
        x_40 : in STD_LOGIC_VECTOR(15 downto 0);
        x_41 : in STD_LOGIC_VECTOR(15 downto 0);
        x_42 : in STD_LOGIC_VECTOR(15 downto 0);
        x_43 : in STD_LOGIC_VECTOR(15 downto 0);
        x_44 : in STD_LOGIC_VECTOR(15 downto 0);
        x_45 : in STD_LOGIC_VECTOR(15 downto 0);
        x_46 : in STD_LOGIC_VECTOR(15 downto 0);
        x_47 : in STD_LOGIC_VECTOR(15 downto 0);
        x_48 : in STD_LOGIC_VECTOR(15 downto 0);
        x_49 : in STD_LOGIC_VECTOR(15 downto 0);
        x_50 : in STD_LOGIC_VECTOR(15 downto 0);
        x_51 : in STD_LOGIC_VECTOR(15 downto 0);
        x_52 : in STD_LOGIC_VECTOR(15 downto 0);
        x_53 : in STD_LOGIC_VECTOR(15 downto 0);
        x_54 : in STD_LOGIC_VECTOR(15 downto 0);
        x_55 : in STD_LOGIC_VECTOR(15 downto 0);
        x_56 : in STD_LOGIC_VECTOR(15 downto 0);
        x_57 : in STD_LOGIC_VECTOR(15 downto 0);
        x_58 : in STD_LOGIC_VECTOR(15 downto 0);
        x_59 : in STD_LOGIC_VECTOR(15 downto 0);
        x_60 : in STD_LOGIC_VECTOR(15 downto 0);
        x_61 : in STD_LOGIC_VECTOR(15 downto 0);
        x_62 : in STD_LOGIC_VECTOR(15 downto 0);
        x_63 : in STD_LOGIC_VECTOR(15 downto 0);
        x_64 : in STD_LOGIC_VECTOR(15 downto 0);
        x_65 : in STD_LOGIC_VECTOR(15 downto 0);
        x_66 : in STD_LOGIC_VECTOR(15 downto 0);
        x_67 : in STD_LOGIC_VECTOR(15 downto 0);
        x_68 : in STD_LOGIC_VECTOR(15 downto 0);
        x_69 : in STD_LOGIC_VECTOR(15 downto 0);
        x_70 : in STD_LOGIC_VECTOR(15 downto 0);
        x_71 : in STD_LOGIC_VECTOR(15 downto 0);
        x_72 : in STD_LOGIC_VECTOR(15 downto 0);
        x_73 : in STD_LOGIC_VECTOR(15 downto 0);
        x_74 : in STD_LOGIC_VECTOR(15 downto 0);
        x_75 : in STD_LOGIC_VECTOR(15 downto 0);
        x_76 : in STD_LOGIC_VECTOR(15 downto 0);
        x_77 : in STD_LOGIC_VECTOR(15 downto 0);
        x_78 : in STD_LOGIC_VECTOR(15 downto 0);
        x_79 : in STD_LOGIC_VECTOR(15 downto 0);
        x_80 : in STD_LOGIC_VECTOR(15 downto 0);
        x_81 : in STD_LOGIC_VECTOR(15 downto 0);
        x_82 : in STD_LOGIC_VECTOR(15 downto 0);
        x_83 : in STD_LOGIC_VECTOR(15 downto 0);
        x_84 : in STD_LOGIC_VECTOR(15 downto 0);
        x_85 : in STD_LOGIC_VECTOR(15 downto 0);
        x_86 : in STD_LOGIC_VECTOR(15 downto 0);
        x_87 : in STD_LOGIC_VECTOR(15 downto 0);
        x_88 : in STD_LOGIC_VECTOR(15 downto 0);
        x_89 : in STD_LOGIC_VECTOR(15 downto 0);
        x_90 : in STD_LOGIC_VECTOR(15 downto 0);
        x_91 : in STD_LOGIC_VECTOR(15 downto 0);
        x_92 : in STD_LOGIC_VECTOR(15 downto 0);
        x_93 : in STD_LOGIC_VECTOR(15 downto 0);
        x_94 : in STD_LOGIC_VECTOR(15 downto 0);
        x_95 : in STD_LOGIC_VECTOR(15 downto 0);
        x_96 : in STD_LOGIC_VECTOR(15 downto 0);
        x_97 : in STD_LOGIC_VECTOR(15 downto 0);
        x_98 : in STD_LOGIC_VECTOR(15 downto 0);
        x_99 : in STD_LOGIC_VECTOR(15 downto 0);
        x_100 : in STD_LOGIC_VECTOR(15 downto 0);
        x_101 : in STD_LOGIC_VECTOR(15 downto 0);
        x_102 : in STD_LOGIC_VECTOR(15 downto 0);
        x_103 : in STD_LOGIC_VECTOR(15 downto 0);
        x_104 : in STD_LOGIC_VECTOR(15 downto 0);
        x_105 : in STD_LOGIC_VECTOR(15 downto 0);
        x_106 : in STD_LOGIC_VECTOR(15 downto 0);
        x_107 : in STD_LOGIC_VECTOR(15 downto 0);
        x_108 : in STD_LOGIC_VECTOR(15 downto 0);
        x_109 : in STD_LOGIC_VECTOR(15 downto 0);
        x_110 : in STD_LOGIC_VECTOR(15 downto 0);
        x_111 : in STD_LOGIC_VECTOR(15 downto 0);
        x_112 : in STD_LOGIC_VECTOR(15 downto 0);
        x_113 : in STD_LOGIC_VECTOR(15 downto 0);
        x_114 : in STD_LOGIC_VECTOR(15 downto 0);
        x_115 : in STD_LOGIC_VECTOR(15 downto 0);
        x_116 : in STD_LOGIC_VECTOR(15 downto 0);
        x_117 : in STD_LOGIC_VECTOR(15 downto 0);
        x_118 : in STD_LOGIC_VECTOR(15 downto 0);
        x_119 : in STD_LOGIC_VECTOR(15 downto 0);
        x_120 : in STD_LOGIC_VECTOR(15 downto 0);
        x_121 : in STD_LOGIC_VECTOR(15 downto 0);
        x_122 : in STD_LOGIC_VECTOR(15 downto 0);
        x_123 : in STD_LOGIC_VECTOR(15 downto 0);
        x_124 : in STD_LOGIC_VECTOR(15 downto 0);
        x_125 : in STD_LOGIC_VECTOR(15 downto 0);
        x_126 : in STD_LOGIC_VECTOR(15 downto 0);
        x_127 : in STD_LOGIC_VECTOR(15 downto 0);
        x_128 : in STD_LOGIC_VECTOR(15 downto 0);
        x_129 : in STD_LOGIC_VECTOR(15 downto 0);
        x_130 : in STD_LOGIC_VECTOR(15 downto 0);
        x_131 : in STD_LOGIC_VECTOR(15 downto 0);
        x_132 : in STD_LOGIC_VECTOR(15 downto 0);
        x_133 : in STD_LOGIC_VECTOR(15 downto 0);
        x_134 : in STD_LOGIC_VECTOR(15 downto 0);
        x_135 : in STD_LOGIC_VECTOR(15 downto 0);
        x_136 : in STD_LOGIC_VECTOR(15 downto 0);
        x_137 : in STD_LOGIC_VECTOR(15 downto 0);
        x_138 : in STD_LOGIC_VECTOR(15 downto 0);
        x_139 : in STD_LOGIC_VECTOR(15 downto 0);
        x_140 : in STD_LOGIC_VECTOR(15 downto 0);
        x_141 : in STD_LOGIC_VECTOR(15 downto 0);
        x_142 : in STD_LOGIC_VECTOR(15 downto 0);
        x_143 : in STD_LOGIC_VECTOR(15 downto 0);
        x_144 : in STD_LOGIC_VECTOR(15 downto 0);
        x_145 : in STD_LOGIC_VECTOR(15 downto 0);
        x_146 : in STD_LOGIC_VECTOR(15 downto 0);
        x_147 : in STD_LOGIC_VECTOR(15 downto 0);
        x_148 : in STD_LOGIC_VECTOR(15 downto 0);
        x_149 : in STD_LOGIC_VECTOR(15 downto 0);
        x_150 : in STD_LOGIC_VECTOR(15 downto 0);
        x_151 : in STD_LOGIC_VECTOR(15 downto 0);
        x_152 : in STD_LOGIC_VECTOR(15 downto 0);
        x_153 : in STD_LOGIC_VECTOR(15 downto 0);
        x_154 : in STD_LOGIC_VECTOR(15 downto 0);
        x_155 : in STD_LOGIC_VECTOR(15 downto 0);
        x_156 : in STD_LOGIC_VECTOR(15 downto 0);
        x_157 : in STD_LOGIC_VECTOR(15 downto 0);
        x_158 : in STD_LOGIC_VECTOR(15 downto 0);
        x_159 : in STD_LOGIC_VECTOR(15 downto 0);
        x_160 : in STD_LOGIC_VECTOR(15 downto 0);
        x_161 : in STD_LOGIC_VECTOR(15 downto 0);
        x_162 : in STD_LOGIC_VECTOR(15 downto 0);
        x_163 : in STD_LOGIC_VECTOR(15 downto 0);
        x_164 : in STD_LOGIC_VECTOR(15 downto 0);
        x_165 : in STD_LOGIC_VECTOR(15 downto 0);
        x_166 : in STD_LOGIC_VECTOR(15 downto 0);
        x_167 : in STD_LOGIC_VECTOR(15 downto 0);
        x_168 : in STD_LOGIC_VECTOR(15 downto 0);
        x_169 : in STD_LOGIC_VECTOR(15 downto 0);
        x_170 : in STD_LOGIC_VECTOR(15 downto 0);
        x_171 : in STD_LOGIC_VECTOR(15 downto 0);
        x_172 : in STD_LOGIC_VECTOR(15 downto 0);
        x_173 : in STD_LOGIC_VECTOR(15 downto 0);
        x_174 : in STD_LOGIC_VECTOR(15 downto 0);
        x_175 : in STD_LOGIC_VECTOR(15 downto 0);
        x_176 : in STD_LOGIC_VECTOR(15 downto 0);
        x_177 : in STD_LOGIC_VECTOR(15 downto 0);
        x_178 : in STD_LOGIC_VECTOR(15 downto 0);
        x_179 : in STD_LOGIC_VECTOR(15 downto 0);
        x_180 : in STD_LOGIC_VECTOR(15 downto 0);
        x_181 : in STD_LOGIC_VECTOR(15 downto 0);
        x_182 : in STD_LOGIC_VECTOR(15 downto 0);
        x_183 : in STD_LOGIC_VECTOR(15 downto 0);
        x_184 : in STD_LOGIC_VECTOR(15 downto 0);
        x_185 : in STD_LOGIC_VECTOR(15 downto 0);
        x_186 : in STD_LOGIC_VECTOR(15 downto 0);
        x_187 : in STD_LOGIC_VECTOR(15 downto 0);
        x_188 : in STD_LOGIC_VECTOR(15 downto 0);
        x_189 : in STD_LOGIC_VECTOR(15 downto 0);
        x_190 : in STD_LOGIC_VECTOR(15 downto 0);
        x_191 : in STD_LOGIC_VECTOR(15 downto 0);
        x_192 : in STD_LOGIC_VECTOR(15 downto 0);
        x_193 : in STD_LOGIC_VECTOR(15 downto 0);
        x_194 : in STD_LOGIC_VECTOR(15 downto 0);
        x_195 : in STD_LOGIC_VECTOR(15 downto 0);
        x_196 : in STD_LOGIC_VECTOR(15 downto 0);
        x_197 : in STD_LOGIC_VECTOR(15 downto 0);
        x_198 : in STD_LOGIC_VECTOR(15 downto 0);
        x_199 : in STD_LOGIC_VECTOR(15 downto 0);
        x_200 : in STD_LOGIC_VECTOR(15 downto 0);
        x_201 : in STD_LOGIC_VECTOR(15 downto 0);
        x_202 : in STD_LOGIC_VECTOR(15 downto 0);
        x_203 : in STD_LOGIC_VECTOR(15 downto 0);
        x_204 : in STD_LOGIC_VECTOR(15 downto 0);
        x_205 : in STD_LOGIC_VECTOR(15 downto 0);
        x_206 : in STD_LOGIC_VECTOR(15 downto 0);
        x_207 : in STD_LOGIC_VECTOR(15 downto 0);
        x_208 : in STD_LOGIC_VECTOR(15 downto 0);
        x_209 : in STD_LOGIC_VECTOR(15 downto 0);
        x_210 : in STD_LOGIC_VECTOR(15 downto 0);
        x_211 : in STD_LOGIC_VECTOR(15 downto 0);
        x_212 : in STD_LOGIC_VECTOR(15 downto 0);
        x_213 : in STD_LOGIC_VECTOR(15 downto 0);
        x_214 : in STD_LOGIC_VECTOR(15 downto 0);
        x_215 : in STD_LOGIC_VECTOR(15 downto 0);
        x_216 : in STD_LOGIC_VECTOR(15 downto 0);
        x_217 : in STD_LOGIC_VECTOR(15 downto 0);
        x_218 : in STD_LOGIC_VECTOR(15 downto 0);
        x_219 : in STD_LOGIC_VECTOR(15 downto 0);
        x_220 : in STD_LOGIC_VECTOR(15 downto 0);
        x_221 : in STD_LOGIC_VECTOR(15 downto 0);
        x_222 : in STD_LOGIC_VECTOR(15 downto 0);
        x_223 : in STD_LOGIC_VECTOR(15 downto 0);
        x_224 : in STD_LOGIC_VECTOR(15 downto 0);
        x_225 : in STD_LOGIC_VECTOR(15 downto 0);
        x_226 : in STD_LOGIC_VECTOR(15 downto 0);
        x_227 : in STD_LOGIC_VECTOR(15 downto 0);
        x_228 : in STD_LOGIC_VECTOR(15 downto 0);
        x_229 : in STD_LOGIC_VECTOR(15 downto 0);
        x_230 : in STD_LOGIC_VECTOR(15 downto 0);
        x_231 : in STD_LOGIC_VECTOR(15 downto 0);
        x_232 : in STD_LOGIC_VECTOR(15 downto 0);
        x_233 : in STD_LOGIC_VECTOR(15 downto 0);
        x_234 : in STD_LOGIC_VECTOR(15 downto 0);
        x_235 : in STD_LOGIC_VECTOR(15 downto 0);
        x_236 : in STD_LOGIC_VECTOR(15 downto 0);
        x_237 : in STD_LOGIC_VECTOR(15 downto 0);
        x_238 : in STD_LOGIC_VECTOR(15 downto 0);
        x_239 : in STD_LOGIC_VECTOR(15 downto 0);
        x_240 : in STD_LOGIC_VECTOR(15 downto 0);
        x_241 : in STD_LOGIC_VECTOR(15 downto 0);
        x_242 : in STD_LOGIC_VECTOR(15 downto 0);
        x_243 : in STD_LOGIC_VECTOR(15 downto 0);
        x_244 : in STD_LOGIC_VECTOR(15 downto 0);
        x_245 : in STD_LOGIC_VECTOR(15 downto 0);
        x_246 : in STD_LOGIC_VECTOR(15 downto 0);
        x_247 : in STD_LOGIC_VECTOR(15 downto 0);
        x_248 : in STD_LOGIC_VECTOR(15 downto 0);
        x_249 : in STD_LOGIC_VECTOR(15 downto 0);
        x_250 : in STD_LOGIC_VECTOR(15 downto 0);
        x_251 : in STD_LOGIC_VECTOR(15 downto 0);
        x_252 : in STD_LOGIC_VECTOR(15 downto 0);
        x_253 : in STD_LOGIC_VECTOR(15 downto 0);
        x_254 : in STD_LOGIC_VECTOR(15 downto 0);
        x_255 : in STD_LOGIC_VECTOR(15 downto 0);
        x_256 : in STD_LOGIC_VECTOR(15 downto 0);
        x_257 : in STD_LOGIC_VECTOR(15 downto 0);
        x_258 : in STD_LOGIC_VECTOR(15 downto 0);
        x_259 : in STD_LOGIC_VECTOR(15 downto 0);
        x_260 : in STD_LOGIC_VECTOR(15 downto 0);
        x_261 : in STD_LOGIC_VECTOR(15 downto 0);
        x_262 : in STD_LOGIC_VECTOR(15 downto 0);
        x_263 : in STD_LOGIC_VECTOR(15 downto 0);
        x_264 : in STD_LOGIC_VECTOR(15 downto 0);
        x_265 : in STD_LOGIC_VECTOR(15 downto 0);
        x_266 : in STD_LOGIC_VECTOR(15 downto 0);
        x_267 : in STD_LOGIC_VECTOR(15 downto 0);
        x_268 : in STD_LOGIC_VECTOR(15 downto 0);
        x_269 : in STD_LOGIC_VECTOR(15 downto 0);
        x_270 : in STD_LOGIC_VECTOR(15 downto 0);
        x_271 : in STD_LOGIC_VECTOR(15 downto 0);
        x_272 : in STD_LOGIC_VECTOR(15 downto 0);
        x_273 : in STD_LOGIC_VECTOR(15 downto 0);
        x_274 : in STD_LOGIC_VECTOR(15 downto 0);
        x_275 : in STD_LOGIC_VECTOR(15 downto 0);
        x_276 : in STD_LOGIC_VECTOR(15 downto 0);
        x_277 : in STD_LOGIC_VECTOR(15 downto 0);
        x_278 : in STD_LOGIC_VECTOR(15 downto 0);
        x_279 : in STD_LOGIC_VECTOR(15 downto 0);
        x_280 : in STD_LOGIC_VECTOR(15 downto 0);
        x_281 : in STD_LOGIC_VECTOR(15 downto 0);
        x_282 : in STD_LOGIC_VECTOR(15 downto 0);
        x_283 : in STD_LOGIC_VECTOR(15 downto 0);
        x_284 : in STD_LOGIC_VECTOR(15 downto 0);
        x_285 : in STD_LOGIC_VECTOR(15 downto 0);
        x_286 : in STD_LOGIC_VECTOR(15 downto 0);
        x_287 : in STD_LOGIC_VECTOR(15 downto 0);
        x_288 : in STD_LOGIC_VECTOR(15 downto 0);
        x_289 : in STD_LOGIC_VECTOR(15 downto 0);
        x_290 : in STD_LOGIC_VECTOR(15 downto 0);
        x_291 : in STD_LOGIC_VECTOR(15 downto 0);
        x_292 : in STD_LOGIC_VECTOR(15 downto 0);
        x_293 : in STD_LOGIC_VECTOR(15 downto 0);
        x_294 : in STD_LOGIC_VECTOR(15 downto 0);
        x_295 : in STD_LOGIC_VECTOR(15 downto 0);
        x_296 : in STD_LOGIC_VECTOR(15 downto 0);
        x_297 : in STD_LOGIC_VECTOR(15 downto 0);
        x_298 : in STD_LOGIC_VECTOR(15 downto 0);
        x_299 : in STD_LOGIC_VECTOR(15 downto 0);
        x_300 : in STD_LOGIC_VECTOR(15 downto 0);
        x_301 : in STD_LOGIC_VECTOR(15 downto 0);
        x_302 : in STD_LOGIC_VECTOR(15 downto 0);
        x_303 : in STD_LOGIC_VECTOR(15 downto 0);
        x_304 : in STD_LOGIC_VECTOR(15 downto 0);
        x_305 : in STD_LOGIC_VECTOR(15 downto 0);
        x_306 : in STD_LOGIC_VECTOR(15 downto 0);
        x_307 : in STD_LOGIC_VECTOR(15 downto 0);
        x_308 : in STD_LOGIC_VECTOR(15 downto 0);
        x_309 : in STD_LOGIC_VECTOR(15 downto 0);
        x_310 : in STD_LOGIC_VECTOR(15 downto 0);
        x_311 : in STD_LOGIC_VECTOR(15 downto 0);
        x_312 : in STD_LOGIC_VECTOR(15 downto 0);
        x_313 : in STD_LOGIC_VECTOR(15 downto 0);
        x_314 : in STD_LOGIC_VECTOR(15 downto 0);
        x_315 : in STD_LOGIC_VECTOR(15 downto 0);
        x_316 : in STD_LOGIC_VECTOR(15 downto 0);
        x_317 : in STD_LOGIC_VECTOR(15 downto 0);
        x_318 : in STD_LOGIC_VECTOR(15 downto 0);
        x_319 : in STD_LOGIC_VECTOR(15 downto 0);
        x_320 : in STD_LOGIC_VECTOR(15 downto 0);
        x_321 : in STD_LOGIC_VECTOR(15 downto 0);
        x_322 : in STD_LOGIC_VECTOR(15 downto 0);
        x_323 : in STD_LOGIC_VECTOR(15 downto 0);
        x_324 : in STD_LOGIC_VECTOR(15 downto 0);
        x_325 : in STD_LOGIC_VECTOR(15 downto 0);
        x_326 : in STD_LOGIC_VECTOR(15 downto 0);
        x_327 : in STD_LOGIC_VECTOR(15 downto 0);
        x_328 : in STD_LOGIC_VECTOR(15 downto 0);
        x_329 : in STD_LOGIC_VECTOR(15 downto 0);
        x_330 : in STD_LOGIC_VECTOR(15 downto 0);
        x_331 : in STD_LOGIC_VECTOR(15 downto 0);
        x_332 : in STD_LOGIC_VECTOR(15 downto 0);
        x_333 : in STD_LOGIC_VECTOR(15 downto 0);
        x_334 : in STD_LOGIC_VECTOR(15 downto 0);
        x_335 : in STD_LOGIC_VECTOR(15 downto 0);
        x_336 : in STD_LOGIC_VECTOR(15 downto 0);
        x_337 : in STD_LOGIC_VECTOR(15 downto 0);
        x_338 : in STD_LOGIC_VECTOR(15 downto 0);
        x_339 : in STD_LOGIC_VECTOR(15 downto 0);
        x_340 : in STD_LOGIC_VECTOR(15 downto 0);
        x_341 : in STD_LOGIC_VECTOR(15 downto 0);
        x_342 : in STD_LOGIC_VECTOR(15 downto 0);
        x_343 : in STD_LOGIC_VECTOR(15 downto 0);
        x_344 : in STD_LOGIC_VECTOR(15 downto 0);
        x_345 : in STD_LOGIC_VECTOR(15 downto 0);
        x_346 : in STD_LOGIC_VECTOR(15 downto 0);
        x_347 : in STD_LOGIC_VECTOR(15 downto 0);
        x_348 : in STD_LOGIC_VECTOR(15 downto 0);
        x_349 : in STD_LOGIC_VECTOR(15 downto 0);
        x_350 : in STD_LOGIC_VECTOR(15 downto 0);
        x_351 : in STD_LOGIC_VECTOR(15 downto 0);
        x_352 : in STD_LOGIC_VECTOR(15 downto 0);
        x_353 : in STD_LOGIC_VECTOR(15 downto 0);
        x_354 : in STD_LOGIC_VECTOR(15 downto 0);
        x_355 : in STD_LOGIC_VECTOR(15 downto 0);
        x_356 : in STD_LOGIC_VECTOR(15 downto 0);
        x_357 : in STD_LOGIC_VECTOR(15 downto 0);
        x_358 : in STD_LOGIC_VECTOR(15 downto 0);
        x_359 : in STD_LOGIC_VECTOR(15 downto 0);
        x_360 : in STD_LOGIC_VECTOR(15 downto 0);
        x_361 : in STD_LOGIC_VECTOR(15 downto 0);
        x_362 : in STD_LOGIC_VECTOR(15 downto 0);
        x_363 : in STD_LOGIC_VECTOR(15 downto 0);
        x_364 : in STD_LOGIC_VECTOR(15 downto 0);
        x_365 : in STD_LOGIC_VECTOR(15 downto 0);
        x_366 : in STD_LOGIC_VECTOR(15 downto 0);
        x_367 : in STD_LOGIC_VECTOR(15 downto 0);
        x_368 : in STD_LOGIC_VECTOR(15 downto 0);
        x_369 : in STD_LOGIC_VECTOR(15 downto 0);
        x_370 : in STD_LOGIC_VECTOR(15 downto 0);
        x_371 : in STD_LOGIC_VECTOR(15 downto 0);
        x_372 : in STD_LOGIC_VECTOR(15 downto 0);
        x_373 : in STD_LOGIC_VECTOR(15 downto 0);
        x_374 : in STD_LOGIC_VECTOR(15 downto 0);
        x_375 : in STD_LOGIC_VECTOR(15 downto 0);
        x_376 : in STD_LOGIC_VECTOR(15 downto 0);
        x_377 : in STD_LOGIC_VECTOR(15 downto 0);
        x_378 : in STD_LOGIC_VECTOR(15 downto 0);
        x_379 : in STD_LOGIC_VECTOR(15 downto 0);
        x_380 : in STD_LOGIC_VECTOR(15 downto 0);
        x_381 : in STD_LOGIC_VECTOR(15 downto 0);
        x_382 : in STD_LOGIC_VECTOR(15 downto 0);
        x_383 : in STD_LOGIC_VECTOR(15 downto 0);
        x_384 : in STD_LOGIC_VECTOR(15 downto 0);
        x_385 : in STD_LOGIC_VECTOR(15 downto 0);
        x_386 : in STD_LOGIC_VECTOR(15 downto 0);
        x_387 : in STD_LOGIC_VECTOR(15 downto 0);
        x_388 : in STD_LOGIC_VECTOR(15 downto 0);
        x_389 : in STD_LOGIC_VECTOR(15 downto 0);
        x_390 : in STD_LOGIC_VECTOR(15 downto 0);
        x_391 : in STD_LOGIC_VECTOR(15 downto 0);
        x_392 : in STD_LOGIC_VECTOR(15 downto 0);
        x_393 : in STD_LOGIC_VECTOR(15 downto 0);
        x_394 : in STD_LOGIC_VECTOR(15 downto 0);
        x_395 : in STD_LOGIC_VECTOR(15 downto 0);
        x_396 : in STD_LOGIC_VECTOR(15 downto 0);
        x_397 : in STD_LOGIC_VECTOR(15 downto 0);
        x_398 : in STD_LOGIC_VECTOR(15 downto 0);
        x_399 : in STD_LOGIC_VECTOR(15 downto 0);
        x_400 : in STD_LOGIC_VECTOR(15 downto 0);
        x_401 : in STD_LOGIC_VECTOR(15 downto 0);
        x_402 : in STD_LOGIC_VECTOR(15 downto 0);
        x_403 : in STD_LOGIC_VECTOR(15 downto 0);
        x_404 : in STD_LOGIC_VECTOR(15 downto 0);
        x_405 : in STD_LOGIC_VECTOR(15 downto 0);
        x_406 : in STD_LOGIC_VECTOR(15 downto 0);
        x_407 : in STD_LOGIC_VECTOR(15 downto 0);
        x_408 : in STD_LOGIC_VECTOR(15 downto 0);
        x_409 : in STD_LOGIC_VECTOR(15 downto 0);
        x_410 : in STD_LOGIC_VECTOR(15 downto 0);
        x_411 : in STD_LOGIC_VECTOR(15 downto 0);
        x_412 : in STD_LOGIC_VECTOR(15 downto 0);
        x_413 : in STD_LOGIC_VECTOR(15 downto 0);
        x_414 : in STD_LOGIC_VECTOR(15 downto 0);
        x_415 : in STD_LOGIC_VECTOR(15 downto 0);
        x_416 : in STD_LOGIC_VECTOR(15 downto 0);
        x_417 : in STD_LOGIC_VECTOR(15 downto 0);
        x_418 : in STD_LOGIC_VECTOR(15 downto 0);
        x_419 : in STD_LOGIC_VECTOR(15 downto 0);
        x_420 : in STD_LOGIC_VECTOR(15 downto 0);
        x_421 : in STD_LOGIC_VECTOR(15 downto 0);
        x_422 : in STD_LOGIC_VECTOR(15 downto 0);
        x_423 : in STD_LOGIC_VECTOR(15 downto 0);
        x_424 : in STD_LOGIC_VECTOR(15 downto 0);
        x_425 : in STD_LOGIC_VECTOR(15 downto 0);
        x_426 : in STD_LOGIC_VECTOR(15 downto 0);
        x_427 : in STD_LOGIC_VECTOR(15 downto 0);
        x_428 : in STD_LOGIC_VECTOR(15 downto 0);
        x_429 : in STD_LOGIC_VECTOR(15 downto 0);
        x_430 : in STD_LOGIC_VECTOR(15 downto 0);
        x_431 : in STD_LOGIC_VECTOR(15 downto 0);
        x_432 : in STD_LOGIC_VECTOR(15 downto 0);
        x_433 : in STD_LOGIC_VECTOR(15 downto 0);
        x_434 : in STD_LOGIC_VECTOR(15 downto 0);
        x_435 : in STD_LOGIC_VECTOR(15 downto 0);
        x_436 : in STD_LOGIC_VECTOR(15 downto 0);
        x_437 : in STD_LOGIC_VECTOR(15 downto 0);
        x_438 : in STD_LOGIC_VECTOR(15 downto 0);
        x_439 : in STD_LOGIC_VECTOR(15 downto 0);
        x_440 : in STD_LOGIC_VECTOR(15 downto 0);
        x_441 : in STD_LOGIC_VECTOR(15 downto 0);
        x_442 : in STD_LOGIC_VECTOR(15 downto 0);
        x_443 : in STD_LOGIC_VECTOR(15 downto 0);
        x_444 : in STD_LOGIC_VECTOR(15 downto 0);
        x_445 : in STD_LOGIC_VECTOR(15 downto 0);
        x_446 : in STD_LOGIC_VECTOR(15 downto 0);
        x_447 : in STD_LOGIC_VECTOR(15 downto 0);
        x_448 : in STD_LOGIC_VECTOR(15 downto 0);
        x_449 : in STD_LOGIC_VECTOR(15 downto 0);
        x_450 : in STD_LOGIC_VECTOR(15 downto 0);
        x_451 : in STD_LOGIC_VECTOR(15 downto 0);
        x_452 : in STD_LOGIC_VECTOR(15 downto 0);
        x_453 : in STD_LOGIC_VECTOR(15 downto 0);
        x_454 : in STD_LOGIC_VECTOR(15 downto 0);
        x_455 : in STD_LOGIC_VECTOR(15 downto 0);
        x_456 : in STD_LOGIC_VECTOR(15 downto 0);
        x_457 : in STD_LOGIC_VECTOR(15 downto 0);
        x_458 : in STD_LOGIC_VECTOR(15 downto 0);
        x_459 : in STD_LOGIC_VECTOR(15 downto 0);
        x_460 : in STD_LOGIC_VECTOR(15 downto 0);
        x_461 : in STD_LOGIC_VECTOR(15 downto 0);
        x_462 : in STD_LOGIC_VECTOR(15 downto 0);
        x_463 : in STD_LOGIC_VECTOR(15 downto 0);
        x_464 : in STD_LOGIC_VECTOR(15 downto 0);
        x_465 : in STD_LOGIC_VECTOR(15 downto 0);
        x_466 : in STD_LOGIC_VECTOR(15 downto 0);
        x_467 : in STD_LOGIC_VECTOR(15 downto 0);
        x_468 : in STD_LOGIC_VECTOR(15 downto 0);
        x_469 : in STD_LOGIC_VECTOR(15 downto 0);
        x_470 : in STD_LOGIC_VECTOR(15 downto 0);
        x_471 : in STD_LOGIC_VECTOR(15 downto 0);
        x_472 : in STD_LOGIC_VECTOR(15 downto 0);
        x_473 : in STD_LOGIC_VECTOR(15 downto 0);
        x_474 : in STD_LOGIC_VECTOR(15 downto 0);
        x_475 : in STD_LOGIC_VECTOR(15 downto 0);
        x_476 : in STD_LOGIC_VECTOR(15 downto 0);
        x_477 : in STD_LOGIC_VECTOR(15 downto 0);
        x_478 : in STD_LOGIC_VECTOR(15 downto 0);
        x_479 : in STD_LOGIC_VECTOR(15 downto 0);
        x_480 : in STD_LOGIC_VECTOR(15 downto 0);
        x_481 : in STD_LOGIC_VECTOR(15 downto 0);
        x_482 : in STD_LOGIC_VECTOR(15 downto 0);
        x_483 : in STD_LOGIC_VECTOR(15 downto 0);
        x_484 : in STD_LOGIC_VECTOR(15 downto 0);
        x_485 : in STD_LOGIC_VECTOR(15 downto 0);
        x_486 : in STD_LOGIC_VECTOR(15 downto 0);
        x_487 : in STD_LOGIC_VECTOR(15 downto 0);
        x_488 : in STD_LOGIC_VECTOR(15 downto 0);
        x_489 : in STD_LOGIC_VECTOR(15 downto 0);
        x_490 : in STD_LOGIC_VECTOR(15 downto 0);
        x_491 : in STD_LOGIC_VECTOR(15 downto 0);
        x_492 : in STD_LOGIC_VECTOR(15 downto 0);
        x_493 : in STD_LOGIC_VECTOR(15 downto 0);
        x_494 : in STD_LOGIC_VECTOR(15 downto 0);
        x_495 : in STD_LOGIC_VECTOR(15 downto 0);
        x_496 : in STD_LOGIC_VECTOR(15 downto 0);
        x_497 : in STD_LOGIC_VECTOR(15 downto 0);
        x_498 : in STD_LOGIC_VECTOR(15 downto 0);
        x_499 : in STD_LOGIC_VECTOR(15 downto 0);
        x_500 : in STD_LOGIC_VECTOR(15 downto 0);
        x_501 : in STD_LOGIC_VECTOR(15 downto 0);
        x_502 : in STD_LOGIC_VECTOR(15 downto 0);
        x_503 : in STD_LOGIC_VECTOR(15 downto 0);
        x_504 : in STD_LOGIC_VECTOR(15 downto 0);
        x_505 : in STD_LOGIC_VECTOR(15 downto 0);
        x_506 : in STD_LOGIC_VECTOR(15 downto 0);
        x_507 : in STD_LOGIC_VECTOR(15 downto 0);
        x_508 : in STD_LOGIC_VECTOR(15 downto 0);
        x_509 : in STD_LOGIC_VECTOR(15 downto 0);
        x_510 : in STD_LOGIC_VECTOR(15 downto 0);
        x_511 : in STD_LOGIC_VECTOR(15 downto 0);
        x_512 : in STD_LOGIC_VECTOR(15 downto 0);
        x_513 : in STD_LOGIC_VECTOR(15 downto 0);
        x_514 : in STD_LOGIC_VECTOR(15 downto 0);
        x_515 : in STD_LOGIC_VECTOR(15 downto 0);
        x_516 : in STD_LOGIC_VECTOR(15 downto 0);
        x_517 : in STD_LOGIC_VECTOR(15 downto 0);
        x_518 : in STD_LOGIC_VECTOR(15 downto 0);
        x_519 : in STD_LOGIC_VECTOR(15 downto 0);
        x_520 : in STD_LOGIC_VECTOR(15 downto 0);
        x_521 : in STD_LOGIC_VECTOR(15 downto 0);
        x_522 : in STD_LOGIC_VECTOR(15 downto 0);
        x_523 : in STD_LOGIC_VECTOR(15 downto 0);
        x_524 : in STD_LOGIC_VECTOR(15 downto 0);
        x_525 : in STD_LOGIC_VECTOR(15 downto 0);
        x_526 : in STD_LOGIC_VECTOR(15 downto 0);
        x_527 : in STD_LOGIC_VECTOR(15 downto 0);
        x_528 : in STD_LOGIC_VECTOR(15 downto 0);
        x_529 : in STD_LOGIC_VECTOR(15 downto 0);
        x_530 : in STD_LOGIC_VECTOR(15 downto 0);
        x_531 : in STD_LOGIC_VECTOR(15 downto 0);
        x_532 : in STD_LOGIC_VECTOR(15 downto 0);
        x_533 : in STD_LOGIC_VECTOR(15 downto 0);
        x_534 : in STD_LOGIC_VECTOR(15 downto 0);
        x_535 : in STD_LOGIC_VECTOR(15 downto 0);
        x_536 : in STD_LOGIC_VECTOR(15 downto 0);
        x_537 : in STD_LOGIC_VECTOR(15 downto 0);
        x_538 : in STD_LOGIC_VECTOR(15 downto 0);
        x_539 : in STD_LOGIC_VECTOR(15 downto 0);
        x_540 : in STD_LOGIC_VECTOR(15 downto 0);
        x_541 : in STD_LOGIC_VECTOR(15 downto 0);
        x_542 : in STD_LOGIC_VECTOR(15 downto 0);
        x_543 : in STD_LOGIC_VECTOR(15 downto 0);
        x_544 : in STD_LOGIC_VECTOR(15 downto 0);
        x_545 : in STD_LOGIC_VECTOR(15 downto 0);
        x_546 : in STD_LOGIC_VECTOR(15 downto 0);
        x_547 : in STD_LOGIC_VECTOR(15 downto 0);
        x_548 : in STD_LOGIC_VECTOR(15 downto 0);
        x_549 : in STD_LOGIC_VECTOR(15 downto 0);
        x_550 : in STD_LOGIC_VECTOR(15 downto 0);
        x_551 : in STD_LOGIC_VECTOR(15 downto 0);
        x_552 : in STD_LOGIC_VECTOR(15 downto 0);
        x_553 : in STD_LOGIC_VECTOR(15 downto 0);
        x_554 : in STD_LOGIC_VECTOR(15 downto 0);
        x_555 : in STD_LOGIC_VECTOR(15 downto 0);
        x_556 : in STD_LOGIC_VECTOR(15 downto 0);
        x_557 : in STD_LOGIC_VECTOR(15 downto 0);
        x_558 : in STD_LOGIC_VECTOR(15 downto 0);
        x_559 : in STD_LOGIC_VECTOR(15 downto 0);
        x_560 : in STD_LOGIC_VECTOR(15 downto 0);
        x_561 : in STD_LOGIC_VECTOR(15 downto 0);
        x_562 : in STD_LOGIC_VECTOR(15 downto 0);
        x_563 : in STD_LOGIC_VECTOR(15 downto 0);
        x_564 : in STD_LOGIC_VECTOR(15 downto 0);
        x_565 : in STD_LOGIC_VECTOR(15 downto 0);
        x_566 : in STD_LOGIC_VECTOR(15 downto 0);
        x_567 : in STD_LOGIC_VECTOR(15 downto 0);
        x_568 : in STD_LOGIC_VECTOR(15 downto 0);
        x_569 : in STD_LOGIC_VECTOR(15 downto 0);
        x_570 : in STD_LOGIC_VECTOR(15 downto 0);
        x_571 : in STD_LOGIC_VECTOR(15 downto 0);
        x_572 : in STD_LOGIC_VECTOR(15 downto 0);
        x_573 : in STD_LOGIC_VECTOR(15 downto 0);
        x_574 : in STD_LOGIC_VECTOR(15 downto 0);
        x_575 : in STD_LOGIC_VECTOR(15 downto 0);
        x_576 : in STD_LOGIC_VECTOR(15 downto 0);
        x_577 : in STD_LOGIC_VECTOR(15 downto 0);
        x_578 : in STD_LOGIC_VECTOR(15 downto 0);
        x_579 : in STD_LOGIC_VECTOR(15 downto 0);
        x_580 : in STD_LOGIC_VECTOR(15 downto 0);
        x_581 : in STD_LOGIC_VECTOR(15 downto 0);
        x_582 : in STD_LOGIC_VECTOR(15 downto 0);
        x_583 : in STD_LOGIC_VECTOR(15 downto 0);
        x_584 : in STD_LOGIC_VECTOR(15 downto 0);
        x_585 : in STD_LOGIC_VECTOR(15 downto 0);
        x_586 : in STD_LOGIC_VECTOR(15 downto 0);
        x_587 : in STD_LOGIC_VECTOR(15 downto 0);
        x_588 : in STD_LOGIC_VECTOR(15 downto 0);
        x_589 : in STD_LOGIC_VECTOR(15 downto 0);
        x_590 : in STD_LOGIC_VECTOR(15 downto 0);
        x_591 : in STD_LOGIC_VECTOR(15 downto 0);
        x_592 : in STD_LOGIC_VECTOR(15 downto 0);
        x_593 : in STD_LOGIC_VECTOR(15 downto 0);
        x_594 : in STD_LOGIC_VECTOR(15 downto 0);
        x_595 : in STD_LOGIC_VECTOR(15 downto 0);
        x_596 : in STD_LOGIC_VECTOR(15 downto 0);
        x_597 : in STD_LOGIC_VECTOR(15 downto 0);
        x_598 : in STD_LOGIC_VECTOR(15 downto 0);
        x_599 : in STD_LOGIC_VECTOR(15 downto 0);
        x_600 : in STD_LOGIC_VECTOR(15 downto 0);
        x_601 : in STD_LOGIC_VECTOR(15 downto 0);
        x_602 : in STD_LOGIC_VECTOR(15 downto 0);
        x_603 : in STD_LOGIC_VECTOR(15 downto 0);
        x_604 : in STD_LOGIC_VECTOR(15 downto 0);
        x_605 : in STD_LOGIC_VECTOR(15 downto 0);
        x_606 : in STD_LOGIC_VECTOR(15 downto 0);
        x_607 : in STD_LOGIC_VECTOR(15 downto 0);
        x_608 : in STD_LOGIC_VECTOR(15 downto 0);
        x_609 : in STD_LOGIC_VECTOR(15 downto 0);
        x_610 : in STD_LOGIC_VECTOR(15 downto 0);
        x_611 : in STD_LOGIC_VECTOR(15 downto 0);
        x_612 : in STD_LOGIC_VECTOR(15 downto 0);
        x_613 : in STD_LOGIC_VECTOR(15 downto 0);
        x_614 : in STD_LOGIC_VECTOR(15 downto 0);
        x_615 : in STD_LOGIC_VECTOR(15 downto 0);
        x_616 : in STD_LOGIC_VECTOR(15 downto 0);
        x_617 : in STD_LOGIC_VECTOR(15 downto 0);
        x_618 : in STD_LOGIC_VECTOR(15 downto 0);
        x_619 : in STD_LOGIC_VECTOR(15 downto 0);
        x_620 : in STD_LOGIC_VECTOR(15 downto 0);
        x_621 : in STD_LOGIC_VECTOR(15 downto 0);
        x_622 : in STD_LOGIC_VECTOR(15 downto 0);
        x_623 : in STD_LOGIC_VECTOR(15 downto 0);
        x_624 : in STD_LOGIC_VECTOR(15 downto 0);
        x_625 : in STD_LOGIC_VECTOR(15 downto 0);
        x_626 : in STD_LOGIC_VECTOR(15 downto 0);
        x_627 : in STD_LOGIC_VECTOR(15 downto 0);
        x_628 : in STD_LOGIC_VECTOR(15 downto 0);
        x_629 : in STD_LOGIC_VECTOR(15 downto 0);
        x_630 : in STD_LOGIC_VECTOR(15 downto 0);
        x_631 : in STD_LOGIC_VECTOR(15 downto 0);
        x_632 : in STD_LOGIC_VECTOR(15 downto 0);
        x_633 : in STD_LOGIC_VECTOR(15 downto 0);
        x_634 : in STD_LOGIC_VECTOR(15 downto 0);
        x_635 : in STD_LOGIC_VECTOR(15 downto 0);
        x_636 : in STD_LOGIC_VECTOR(15 downto 0);
        x_637 : in STD_LOGIC_VECTOR(15 downto 0);
        x_638 : in STD_LOGIC_VECTOR(15 downto 0);
        x_639 : in STD_LOGIC_VECTOR(15 downto 0);
        x_640 : in STD_LOGIC_VECTOR(15 downto 0);
        x_641 : in STD_LOGIC_VECTOR(15 downto 0);
        x_642 : in STD_LOGIC_VECTOR(15 downto 0);
        x_643 : in STD_LOGIC_VECTOR(15 downto 0);
        x_644 : in STD_LOGIC_VECTOR(15 downto 0);
        x_645 : in STD_LOGIC_VECTOR(15 downto 0);
        x_646 : in STD_LOGIC_VECTOR(15 downto 0);
        x_647 : in STD_LOGIC_VECTOR(15 downto 0);
        x_648 : in STD_LOGIC_VECTOR(15 downto 0);
        x_649 : in STD_LOGIC_VECTOR(15 downto 0);
        x_650 : in STD_LOGIC_VECTOR(15 downto 0);
        x_651 : in STD_LOGIC_VECTOR(15 downto 0);
        x_652 : in STD_LOGIC_VECTOR(15 downto 0);
        x_653 : in STD_LOGIC_VECTOR(15 downto 0);
        x_654 : in STD_LOGIC_VECTOR(15 downto 0);
        x_655 : in STD_LOGIC_VECTOR(15 downto 0);
        x_656 : in STD_LOGIC_VECTOR(15 downto 0);
        x_657 : in STD_LOGIC_VECTOR(15 downto 0);
        x_658 : in STD_LOGIC_VECTOR(15 downto 0);
        x_659 : in STD_LOGIC_VECTOR(15 downto 0);
        x_660 : in STD_LOGIC_VECTOR(15 downto 0);
        x_661 : in STD_LOGIC_VECTOR(15 downto 0);
        x_662 : in STD_LOGIC_VECTOR(15 downto 0);
        x_663 : in STD_LOGIC_VECTOR(15 downto 0);
        x_664 : in STD_LOGIC_VECTOR(15 downto 0);
        x_665 : in STD_LOGIC_VECTOR(15 downto 0);
        x_666 : in STD_LOGIC_VECTOR(15 downto 0);
        x_667 : in STD_LOGIC_VECTOR(15 downto 0);
        x_668 : in STD_LOGIC_VECTOR(15 downto 0);
        x_669 : in STD_LOGIC_VECTOR(15 downto 0);
        x_670 : in STD_LOGIC_VECTOR(15 downto 0);
        x_671 : in STD_LOGIC_VECTOR(15 downto 0);
        x_672 : in STD_LOGIC_VECTOR(15 downto 0);
        x_673 : in STD_LOGIC_VECTOR(15 downto 0);
        x_674 : in STD_LOGIC_VECTOR(15 downto 0);
        x_675 : in STD_LOGIC_VECTOR(15 downto 0);
        x_676 : in STD_LOGIC_VECTOR(15 downto 0);
        x_677 : in STD_LOGIC_VECTOR(15 downto 0);
        x_678 : in STD_LOGIC_VECTOR(15 downto 0);
        x_679 : in STD_LOGIC_VECTOR(15 downto 0);
        x_680 : in STD_LOGIC_VECTOR(15 downto 0);
        x_681 : in STD_LOGIC_VECTOR(15 downto 0);
        x_682 : in STD_LOGIC_VECTOR(15 downto 0);
        x_683 : in STD_LOGIC_VECTOR(15 downto 0);
        x_684 : in STD_LOGIC_VECTOR(15 downto 0);
        x_685 : in STD_LOGIC_VECTOR(15 downto 0);
        x_686 : in STD_LOGIC_VECTOR(15 downto 0);
        x_687 : in STD_LOGIC_VECTOR(15 downto 0);
        x_688 : in STD_LOGIC_VECTOR(15 downto 0);
        x_689 : in STD_LOGIC_VECTOR(15 downto 0);
        x_690 : in STD_LOGIC_VECTOR(15 downto 0);
        x_691 : in STD_LOGIC_VECTOR(15 downto 0);
        x_692 : in STD_LOGIC_VECTOR(15 downto 0);
        x_693 : in STD_LOGIC_VECTOR(15 downto 0);
        x_694 : in STD_LOGIC_VECTOR(15 downto 0);
        x_695 : in STD_LOGIC_VECTOR(15 downto 0);
        x_696 : in STD_LOGIC_VECTOR(15 downto 0);
        x_697 : in STD_LOGIC_VECTOR(15 downto 0);
        x_698 : in STD_LOGIC_VECTOR(15 downto 0);
        x_699 : in STD_LOGIC_VECTOR(15 downto 0);
        x_700 : in STD_LOGIC_VECTOR(15 downto 0);
        x_701 : in STD_LOGIC_VECTOR(15 downto 0);
        x_702 : in STD_LOGIC_VECTOR(15 downto 0);
        x_703 : in STD_LOGIC_VECTOR(15 downto 0);
        x_704 : in STD_LOGIC_VECTOR(15 downto 0);
        x_705 : in STD_LOGIC_VECTOR(15 downto 0);
        x_706 : in STD_LOGIC_VECTOR(15 downto 0);
        x_707 : in STD_LOGIC_VECTOR(15 downto 0);
        x_708 : in STD_LOGIC_VECTOR(15 downto 0);
        x_709 : in STD_LOGIC_VECTOR(15 downto 0);
        x_710 : in STD_LOGIC_VECTOR(15 downto 0);
        x_711 : in STD_LOGIC_VECTOR(15 downto 0);
        x_712 : in STD_LOGIC_VECTOR(15 downto 0);
        x_713 : in STD_LOGIC_VECTOR(15 downto 0);
        x_714 : in STD_LOGIC_VECTOR(15 downto 0);
        x_715 : in STD_LOGIC_VECTOR(15 downto 0);
        x_716 : in STD_LOGIC_VECTOR(15 downto 0);
        x_717 : in STD_LOGIC_VECTOR(15 downto 0);
        x_718 : in STD_LOGIC_VECTOR(15 downto 0);
        x_719 : in STD_LOGIC_VECTOR(15 downto 0);
        x_720 : in STD_LOGIC_VECTOR(15 downto 0);
        x_721 : in STD_LOGIC_VECTOR(15 downto 0);
        x_722 : in STD_LOGIC_VECTOR(15 downto 0);
        x_723 : in STD_LOGIC_VECTOR(15 downto 0);
        x_724 : in STD_LOGIC_VECTOR(15 downto 0);
        x_725 : in STD_LOGIC_VECTOR(15 downto 0);
        x_726 : in STD_LOGIC_VECTOR(15 downto 0);
        x_727 : in STD_LOGIC_VECTOR(15 downto 0);
        x_728 : in STD_LOGIC_VECTOR(15 downto 0);
        x_729 : in STD_LOGIC_VECTOR(15 downto 0);
        x_730 : in STD_LOGIC_VECTOR(15 downto 0);
        x_731 : in STD_LOGIC_VECTOR(15 downto 0);
        x_732 : in STD_LOGIC_VECTOR(15 downto 0);
        x_733 : in STD_LOGIC_VECTOR(15 downto 0);
        x_734 : in STD_LOGIC_VECTOR(15 downto 0);
        x_735 : in STD_LOGIC_VECTOR(15 downto 0);
        x_736 : in STD_LOGIC_VECTOR(15 downto 0);
        x_737 : in STD_LOGIC_VECTOR(15 downto 0);
        x_738 : in STD_LOGIC_VECTOR(15 downto 0);
        x_739 : in STD_LOGIC_VECTOR(15 downto 0);
        x_740 : in STD_LOGIC_VECTOR(15 downto 0);
        x_741 : in STD_LOGIC_VECTOR(15 downto 0);
        x_742 : in STD_LOGIC_VECTOR(15 downto 0);
        x_743 : in STD_LOGIC_VECTOR(15 downto 0);
        x_744 : in STD_LOGIC_VECTOR(15 downto 0);
        x_745 : in STD_LOGIC_VECTOR(15 downto 0);
        x_746 : in STD_LOGIC_VECTOR(15 downto 0);
        x_747 : in STD_LOGIC_VECTOR(15 downto 0);
        x_748 : in STD_LOGIC_VECTOR(15 downto 0);
        x_749 : in STD_LOGIC_VECTOR(15 downto 0);
        x_750 : in STD_LOGIC_VECTOR(15 downto 0);
        x_751 : in STD_LOGIC_VECTOR(15 downto 0);
        x_752 : in STD_LOGIC_VECTOR(15 downto 0);
        x_753 : in STD_LOGIC_VECTOR(15 downto 0);
        x_754 : in STD_LOGIC_VECTOR(15 downto 0);
        x_755 : in STD_LOGIC_VECTOR(15 downto 0);
        x_756 : in STD_LOGIC_VECTOR(15 downto 0);
        x_757 : in STD_LOGIC_VECTOR(15 downto 0);
        x_758 : in STD_LOGIC_VECTOR(15 downto 0);
        x_759 : in STD_LOGIC_VECTOR(15 downto 0);
        x_760 : in STD_LOGIC_VECTOR(15 downto 0);
        x_761 : in STD_LOGIC_VECTOR(15 downto 0);
        x_762 : in STD_LOGIC_VECTOR(15 downto 0);
        x_763 : in STD_LOGIC_VECTOR(15 downto 0);
        x_764 : in STD_LOGIC_VECTOR(15 downto 0);
        x_765 : in STD_LOGIC_VECTOR(15 downto 0);
        x_766 : in STD_LOGIC_VECTOR(15 downto 0);
        x_767 : in STD_LOGIC_VECTOR(15 downto 0);
        x_768 : in STD_LOGIC_VECTOR(15 downto 0);
        x_769 : in STD_LOGIC_VECTOR(15 downto 0);
        x_770 : in STD_LOGIC_VECTOR(15 downto 0);
        x_771 : in STD_LOGIC_VECTOR(15 downto 0);
        x_772 : in STD_LOGIC_VECTOR(15 downto 0);
        x_773 : in STD_LOGIC_VECTOR(15 downto 0);
        x_774 : in STD_LOGIC_VECTOR(15 downto 0);
        x_775 : in STD_LOGIC_VECTOR(15 downto 0);
        x_776 : in STD_LOGIC_VECTOR(15 downto 0);
        x_777 : in STD_LOGIC_VECTOR(15 downto 0);
        x_778 : in STD_LOGIC_VECTOR(15 downto 0);
        x_779 : in STD_LOGIC_VECTOR(15 downto 0);
        x_780 : in STD_LOGIC_VECTOR(15 downto 0);
        x_781 : in STD_LOGIC_VECTOR(15 downto 0);
        x_782 : in STD_LOGIC_VECTOR(15 downto 0);
        x_783 : in STD_LOGIC_VECTOR(15 downto 0);
        y : out STD_LOGIC_VECTOR(3 downto 0));
end component fully_connected_layer;

begin
   ut0_lstm_layer: lstm_layer port map(
       clk=> clk,
       x_0=> x_0,
       x_1=> x_1,
       x_2=> x_2,
       x_3=> x_3,
       x_4=> x_4,
       x_5=> x_5,
       x_6=> x_6,
       x_7=> x_7,
       x_8=> x_8,
       x_9=> x_9,
       x_10=> x_10,
       x_11=> x_11,
       x_12=> x_12,
       x_13=> x_13,
       x_14=> x_14,
       x_15=> x_15,
       x_16=> x_16,
       x_17=> x_17,
       x_18=> x_18,
       x_19=> x_19,
       x_20=> x_20,
       x_21=> x_21,
       x_22=> x_22,
       x_23=> x_23,
       x_24=> x_24,
       x_25=> x_25,
       x_26=> x_26,
       x_27=> x_27,
       x_28=> x_28,
       x_29=> x_29,
       x_30=> x_30,
       x_31=> x_31,
       x_32=> x_32,
       x_33=> x_33,
       x_34=> x_34,
       x_35=> x_35,
       x_36=> x_36,
       x_37=> x_37,
       x_38=> x_38,
       x_39=> x_39,
       x_40=> x_40,
       x_41=> x_41,
       x_42=> x_42,
       x_43=> x_43,
       x_44=> x_44,
       x_45=> x_45,
       x_46=> x_46,
       x_47=> x_47,
       x_48=> x_48,
       x_49=> x_49,
       x_50=> x_50,
       x_51=> x_51,
       x_52=> x_52,
       x_53=> x_53,
       x_54=> x_54,
       x_55=> x_55,
       x_56=> x_56,
       x_57=> x_57,
       x_58=> x_58,
       x_59=> x_59,
       x_60=> x_60,
       x_61=> x_61,
       x_62=> x_62,
       x_63=> x_63,
       x_64=> x_64,
       x_65=> x_65,
       x_66=> x_66,
       x_67=> x_67,
       x_68=> x_68,
       x_69=> x_69,
       x_70=> x_70,
       x_71=> x_71,
       x_72=> x_72,
       x_73=> x_73,
       x_74=> x_74,
       x_75=> x_75,
       x_76=> x_76,
       x_77=> x_77,
       x_78=> x_78,
       x_79=> x_79,
       x_80=> x_80,
       x_81=> x_81,
       x_82=> x_82,
       x_83=> x_83,
       x_84=> x_84,
       x_85=> x_85,
       x_86=> x_86,
       x_87=> x_87,
       x_88=> x_88,
       x_89=> x_89,
       x_90=> x_90,
       x_91=> x_91,
       x_92=> x_92,
       x_93=> x_93,
       x_94=> x_94,
       x_95=> x_95,
       x_96=> x_96,
       x_97=> x_97,
       x_98=> x_98,
       x_99=> x_99,
       x_100=> x_100,
       x_101=> x_101,
       x_102=> x_102,
       x_103=> x_103,
       x_104=> x_104,
       x_105=> x_105,
       x_106=> x_106,
       x_107=> x_107,
       x_108=> x_108,
       x_109=> x_109,
       x_110=> x_110,
       x_111=> x_111,
       x_112=> x_112,
       x_113=> x_113,
       x_114=> x_114,
       x_115=> x_115,
       x_116=> x_116,
       x_117=> x_117,
       x_118=> x_118,
       x_119=> x_119,
       x_120=> x_120,
       x_121=> x_121,
       x_122=> x_122,
       x_123=> x_123,
       x_124=> x_124,
       x_125=> x_125,
       x_126=> x_126,
       x_127=> x_127,
       x_128=> x_128,
       x_129=> x_129,
       x_130=> x_130,
       x_131=> x_131,
       x_132=> x_132,
       x_133=> x_133,
       x_134=> x_134,
       x_135=> x_135,
       x_136=> x_136,
       x_137=> x_137,
       x_138=> x_138,
       x_139=> x_139,
       x_140=> x_140,
       x_141=> x_141,
       x_142=> x_142,
       x_143=> x_143,
       x_144=> x_144,
       x_145=> x_145,
       x_146=> x_146,
       x_147=> x_147,
       x_148=> x_148,
       x_149=> x_149,
       x_150=> x_150,
       x_151=> x_151,
       x_152=> x_152,
       x_153=> x_153,
       x_154=> x_154,
       x_155=> x_155,
       x_156=> x_156,
       x_157=> x_157,
       x_158=> x_158,
       x_159=> x_159,
       x_160=> x_160,
       x_161=> x_161,
       x_162=> x_162,
       x_163=> x_163,
       x_164=> x_164,
       x_165=> x_165,
       x_166=> x_166,
       x_167=> x_167,
       x_168=> x_168,
       x_169=> x_169,
       x_170=> x_170,
       x_171=> x_171,
       x_172=> x_172,
       x_173=> x_173,
       x_174=> x_174,
       x_175=> x_175,
       x_176=> x_176,
       x_177=> x_177,
       x_178=> x_178,
       x_179=> x_179,
       x_180=> x_180,
       x_181=> x_181,
       x_182=> x_182,
       x_183=> x_183,
       x_184=> x_184,
       x_185=> x_185,
       x_186=> x_186,
       x_187=> x_187,
       x_188=> x_188,
       x_189=> x_189,
       x_190=> x_190,
       x_191=> x_191,
       x_192=> x_192,
       x_193=> x_193,
       x_194=> x_194,
       x_195=> x_195,
       x_196=> x_196,
       x_197=> x_197,
       x_198=> x_198,
       x_199=> x_199,
       x_200=> x_200,
       x_201=> x_201,
       x_202=> x_202,
       x_203=> x_203,
       x_204=> x_204,
       x_205=> x_205,
       x_206=> x_206,
       x_207=> x_207,
       x_208=> x_208,
       x_209=> x_209,
       x_210=> x_210,
       x_211=> x_211,
       x_212=> x_212,
       x_213=> x_213,
       x_214=> x_214,
       x_215=> x_215,
       x_216=> x_216,
       x_217=> x_217,
       x_218=> x_218,
       x_219=> x_219,
       x_220=> x_220,
       x_221=> x_221,
       x_222=> x_222,
       x_223=> x_223,
       x_224=> x_224,
       x_225=> x_225,
       x_226=> x_226,
       x_227=> x_227,
       x_228=> x_228,
       x_229=> x_229,
       x_230=> x_230,
       x_231=> x_231,
       x_232=> x_232,
       x_233=> x_233,
       x_234=> x_234,
       x_235=> x_235,
       x_236=> x_236,
       x_237=> x_237,
       x_238=> x_238,
       x_239=> x_239,
       x_240=> x_240,
       x_241=> x_241,
       x_242=> x_242,
       x_243=> x_243,
       x_244=> x_244,
       x_245=> x_245,
       x_246=> x_246,
       x_247=> x_247,
       x_248=> x_248,
       x_249=> x_249,
       x_250=> x_250,
       x_251=> x_251,
       x_252=> x_252,
       x_253=> x_253,
       x_254=> x_254,
       x_255=> x_255,
       x_256=> x_256,
       x_257=> x_257,
       x_258=> x_258,
       x_259=> x_259,
       x_260=> x_260,
       x_261=> x_261,
       x_262=> x_262,
       x_263=> x_263,
       x_264=> x_264,
       x_265=> x_265,
       x_266=> x_266,
       x_267=> x_267,
       x_268=> x_268,
       x_269=> x_269,
       x_270=> x_270,
       x_271=> x_271,
       x_272=> x_272,
       x_273=> x_273,
       x_274=> x_274,
       x_275=> x_275,
       x_276=> x_276,
       x_277=> x_277,
       x_278=> x_278,
       x_279=> x_279,
       x_280=> x_280,
       x_281=> x_281,
       x_282=> x_282,
       x_283=> x_283,
       x_284=> x_284,
       x_285=> x_285,
       x_286=> x_286,
       x_287=> x_287,
       x_288=> x_288,
       x_289=> x_289,
       x_290=> x_290,
       x_291=> x_291,
       x_292=> x_292,
       x_293=> x_293,
       x_294=> x_294,
       x_295=> x_295,
       x_296=> x_296,
       x_297=> x_297,
       x_298=> x_298,
       x_299=> x_299,
       x_300=> x_300,
       x_301=> x_301,
       x_302=> x_302,
       x_303=> x_303,
       x_304=> x_304,
       x_305=> x_305,
       x_306=> x_306,
       x_307=> x_307,
       x_308=> x_308,
       x_309=> x_309,
       x_310=> x_310,
       x_311=> x_311,
       x_312=> x_312,
       x_313=> x_313,
       x_314=> x_314,
       x_315=> x_315,
       x_316=> x_316,
       x_317=> x_317,
       x_318=> x_318,
       x_319=> x_319,
       x_320=> x_320,
       x_321=> x_321,
       x_322=> x_322,
       x_323=> x_323,
       x_324=> x_324,
       x_325=> x_325,
       x_326=> x_326,
       x_327=> x_327,
       x_328=> x_328,
       x_329=> x_329,
       x_330=> x_330,
       x_331=> x_331,
       x_332=> x_332,
       x_333=> x_333,
       x_334=> x_334,
       x_335=> x_335,
       x_336=> x_336,
       x_337=> x_337,
       x_338=> x_338,
       x_339=> x_339,
       x_340=> x_340,
       x_341=> x_341,
       x_342=> x_342,
       x_343=> x_343,
       x_344=> x_344,
       x_345=> x_345,
       x_346=> x_346,
       x_347=> x_347,
       x_348=> x_348,
       x_349=> x_349,
       x_350=> x_350,
       x_351=> x_351,
       x_352=> x_352,
       x_353=> x_353,
       x_354=> x_354,
       x_355=> x_355,
       x_356=> x_356,
       x_357=> x_357,
       x_358=> x_358,
       x_359=> x_359,
       x_360=> x_360,
       x_361=> x_361,
       x_362=> x_362,
       x_363=> x_363,
       x_364=> x_364,
       x_365=> x_365,
       x_366=> x_366,
       x_367=> x_367,
       x_368=> x_368,
       x_369=> x_369,
       x_370=> x_370,
       x_371=> x_371,
       x_372=> x_372,
       x_373=> x_373,
       x_374=> x_374,
       x_375=> x_375,
       x_376=> x_376,
       x_377=> x_377,
       x_378=> x_378,
       x_379=> x_379,
       x_380=> x_380,
       x_381=> x_381,
       x_382=> x_382,
       x_383=> x_383,
       x_384=> x_384,
       x_385=> x_385,
       x_386=> x_386,
       x_387=> x_387,
       x_388=> x_388,
       x_389=> x_389,
       x_390=> x_390,
       x_391=> x_391,
       x_392=> x_392,
       x_393=> x_393,
       x_394=> x_394,
       x_395=> x_395,
       x_396=> x_396,
       x_397=> x_397,
       x_398=> x_398,
       x_399=> x_399,
       x_400=> x_400,
       x_401=> x_401,
       x_402=> x_402,
       x_403=> x_403,
       x_404=> x_404,
       x_405=> x_405,
       x_406=> x_406,
       x_407=> x_407,
       x_408=> x_408,
       x_409=> x_409,
       x_410=> x_410,
       x_411=> x_411,
       x_412=> x_412,
       x_413=> x_413,
       x_414=> x_414,
       x_415=> x_415,
       x_416=> x_416,
       x_417=> x_417,
       x_418=> x_418,
       x_419=> x_419,
       x_420=> x_420,
       x_421=> x_421,
       x_422=> x_422,
       x_423=> x_423,
       x_424=> x_424,
       x_425=> x_425,
       x_426=> x_426,
       x_427=> x_427,
       x_428=> x_428,
       x_429=> x_429,
       x_430=> x_430,
       x_431=> x_431,
       x_432=> x_432,
       x_433=> x_433,
       x_434=> x_434,
       x_435=> x_435,
       x_436=> x_436,
       x_437=> x_437,
       x_438=> x_438,
       x_439=> x_439,
       x_440=> x_440,
       x_441=> x_441,
       x_442=> x_442,
       x_443=> x_443,
       x_444=> x_444,
       x_445=> x_445,
       x_446=> x_446,
       x_447=> x_447,
       x_448=> x_448,
       x_449=> x_449,
       x_450=> x_450,
       x_451=> x_451,
       x_452=> x_452,
       x_453=> x_453,
       x_454=> x_454,
       x_455=> x_455,
       x_456=> x_456,
       x_457=> x_457,
       x_458=> x_458,
       x_459=> x_459,
       x_460=> x_460,
       x_461=> x_461,
       x_462=> x_462,
       x_463=> x_463,
       x_464=> x_464,
       x_465=> x_465,
       x_466=> x_466,
       x_467=> x_467,
       x_468=> x_468,
       x_469=> x_469,
       x_470=> x_470,
       x_471=> x_471,
       x_472=> x_472,
       x_473=> x_473,
       x_474=> x_474,
       x_475=> x_475,
       x_476=> x_476,
       x_477=> x_477,
       x_478=> x_478,
       x_479=> x_479,
       x_480=> x_480,
       x_481=> x_481,
       x_482=> x_482,
       x_483=> x_483,
       x_484=> x_484,
       x_485=> x_485,
       x_486=> x_486,
       x_487=> x_487,
       x_488=> x_488,
       x_489=> x_489,
       x_490=> x_490,
       x_491=> x_491,
       x_492=> x_492,
       x_493=> x_493,
       x_494=> x_494,
       x_495=> x_495,
       x_496=> x_496,
       x_497=> x_497,
       x_498=> x_498,
       x_499=> x_499,
       x_500=> x_500,
       x_501=> x_501,
       x_502=> x_502,
       x_503=> x_503,
       x_504=> x_504,
       x_505=> x_505,
       x_506=> x_506,
       x_507=> x_507,
       x_508=> x_508,
       x_509=> x_509,
       x_510=> x_510,
       x_511=> x_511,
       x_512=> x_512,
       x_513=> x_513,
       x_514=> x_514,
       x_515=> x_515,
       x_516=> x_516,
       x_517=> x_517,
       x_518=> x_518,
       x_519=> x_519,
       x_520=> x_520,
       x_521=> x_521,
       x_522=> x_522,
       x_523=> x_523,
       x_524=> x_524,
       x_525=> x_525,
       x_526=> x_526,
       x_527=> x_527,
       x_528=> x_528,
       x_529=> x_529,
       x_530=> x_530,
       x_531=> x_531,
       x_532=> x_532,
       x_533=> x_533,
       x_534=> x_534,
       x_535=> x_535,
       x_536=> x_536,
       x_537=> x_537,
       x_538=> x_538,
       x_539=> x_539,
       x_540=> x_540,
       x_541=> x_541,
       x_542=> x_542,
       x_543=> x_543,
       x_544=> x_544,
       x_545=> x_545,
       x_546=> x_546,
       x_547=> x_547,
       x_548=> x_548,
       x_549=> x_549,
       x_550=> x_550,
       x_551=> x_551,
       x_552=> x_552,
       x_553=> x_553,
       x_554=> x_554,
       x_555=> x_555,
       x_556=> x_556,
       x_557=> x_557,
       x_558=> x_558,
       x_559=> x_559,
       x_560=> x_560,
       x_561=> x_561,
       x_562=> x_562,
       x_563=> x_563,
       x_564=> x_564,
       x_565=> x_565,
       x_566=> x_566,
       x_567=> x_567,
       x_568=> x_568,
       x_569=> x_569,
       x_570=> x_570,
       x_571=> x_571,
       x_572=> x_572,
       x_573=> x_573,
       x_574=> x_574,
       x_575=> x_575,
       x_576=> x_576,
       x_577=> x_577,
       x_578=> x_578,
       x_579=> x_579,
       x_580=> x_580,
       x_581=> x_581,
       x_582=> x_582,
       x_583=> x_583,
       x_584=> x_584,
       x_585=> x_585,
       x_586=> x_586,
       x_587=> x_587,
       x_588=> x_588,
       x_589=> x_589,
       x_590=> x_590,
       x_591=> x_591,
       x_592=> x_592,
       x_593=> x_593,
       x_594=> x_594,
       x_595=> x_595,
       x_596=> x_596,
       x_597=> x_597,
       x_598=> x_598,
       x_599=> x_599,
       x_600=> x_600,
       x_601=> x_601,
       x_602=> x_602,
       x_603=> x_603,
       x_604=> x_604,
       x_605=> x_605,
       x_606=> x_606,
       x_607=> x_607,
       x_608=> x_608,
       x_609=> x_609,
       x_610=> x_610,
       x_611=> x_611,
       x_612=> x_612,
       x_613=> x_613,
       x_614=> x_614,
       x_615=> x_615,
       x_616=> x_616,
       x_617=> x_617,
       x_618=> x_618,
       x_619=> x_619,
       x_620=> x_620,
       x_621=> x_621,
       x_622=> x_622,
       x_623=> x_623,
       x_624=> x_624,
       x_625=> x_625,
       x_626=> x_626,
       x_627=> x_627,
       x_628=> x_628,
       x_629=> x_629,
       x_630=> x_630,
       x_631=> x_631,
       x_632=> x_632,
       x_633=> x_633,
       x_634=> x_634,
       x_635=> x_635,
       x_636=> x_636,
       x_637=> x_637,
       x_638=> x_638,
       x_639=> x_639,
       x_640=> x_640,
       x_641=> x_641,
       x_642=> x_642,
       x_643=> x_643,
       x_644=> x_644,
       x_645=> x_645,
       x_646=> x_646,
       x_647=> x_647,
       x_648=> x_648,
       x_649=> x_649,
       x_650=> x_650,
       x_651=> x_651,
       x_652=> x_652,
       x_653=> x_653,
       x_654=> x_654,
       x_655=> x_655,
       x_656=> x_656,
       x_657=> x_657,
       x_658=> x_658,
       x_659=> x_659,
       x_660=> x_660,
       x_661=> x_661,
       x_662=> x_662,
       x_663=> x_663,
       x_664=> x_664,
       x_665=> x_665,
       x_666=> x_666,
       x_667=> x_667,
       x_668=> x_668,
       x_669=> x_669,
       x_670=> x_670,
       x_671=> x_671,
       x_672=> x_672,
       x_673=> x_673,
       x_674=> x_674,
       x_675=> x_675,
       x_676=> x_676,
       x_677=> x_677,
       x_678=> x_678,
       x_679=> x_679,
       x_680=> x_680,
       x_681=> x_681,
       x_682=> x_682,
       x_683=> x_683,
       x_684=> x_684,
       x_685=> x_685,
       x_686=> x_686,
       x_687=> x_687,
       x_688=> x_688,
       x_689=> x_689,
       x_690=> x_690,
       x_691=> x_691,
       x_692=> x_692,
       x_693=> x_693,
       x_694=> x_694,
       x_695=> x_695,
       x_696=> x_696,
       x_697=> x_697,
       x_698=> x_698,
       x_699=> x_699,
       x_700=> x_700,
       x_701=> x_701,
       x_702=> x_702,
       x_703=> x_703,
       x_704=> x_704,
       x_705=> x_705,
       x_706=> x_706,
       x_707=> x_707,
       x_708=> x_708,
       x_709=> x_709,
       x_710=> x_710,
       x_711=> x_711,
       x_712=> x_712,
       x_713=> x_713,
       x_714=> x_714,
       x_715=> x_715,
       x_716=> x_716,
       x_717=> x_717,
       x_718=> x_718,
       x_719=> x_719,
       x_720=> x_720,
       x_721=> x_721,
       x_722=> x_722,
       x_723=> x_723,
       x_724=> x_724,
       x_725=> x_725,
       x_726=> x_726,
       x_727=> x_727,
       x_728=> x_728,
       x_729=> x_729,
       x_730=> x_730,
       x_731=> x_731,
       x_732=> x_732,
       x_733=> x_733,
       x_734=> x_734,
       x_735=> x_735,
       x_736=> x_736,
       x_737=> x_737,
       x_738=> x_738,
       x_739=> x_739,
       x_740=> x_740,
       x_741=> x_741,
       x_742=> x_742,
       x_743=> x_743,
       x_744=> x_744,
       x_745=> x_745,
       x_746=> x_746,
       x_747=> x_747,
       x_748=> x_748,
       x_749=> x_749,
       x_750=> x_750,
       x_751=> x_751,
       x_752=> x_752,
       x_753=> x_753,
       x_754=> x_754,
       x_755=> x_755,
       x_756=> x_756,
       x_757=> x_757,
       x_758=> x_758,
       x_759=> x_759,
       x_760=> x_760,
       x_761=> x_761,
       x_762=> x_762,
       x_763=> x_763,
       x_764=> x_764,
       x_765=> x_765,
       x_766=> x_766,
       x_767=> x_767,
       x_768=> x_768,
       x_769=> x_769,
       x_770=> x_770,
       x_771=> x_771,
       x_772=> x_772,
       x_773=> x_773,
       x_774=> x_774,
       x_775=> x_775,
       x_776=> x_776,
       x_777=> x_777,
       x_778=> x_778,
       x_779=> x_779,
       x_780=> x_780,
       x_781=> x_781,
       x_782=> x_782,
       x_783=> x_783,
       y_0=> store_value_0,
       y_1=> store_value_1,
       y_2=> store_value_2,
       y_3=> store_value_3,
       y_4=> store_value_4,
       y_5=> store_value_5,
       y_6=> store_value_6,
       y_7=> store_value_7,
       y_8=> store_value_8,
       y_9=> store_value_9,
       y_10=> store_value_10,
       y_11=> store_value_11,
       y_12=> store_value_12,
       y_13=> store_value_13,
       y_14=> store_value_14,
       y_15=> store_value_15,
       y_16=> store_value_16,
       y_17=> store_value_17,
       y_18=> store_value_18,
       y_19=> store_value_19,
       y_20=> store_value_20,
       y_21=> store_value_21,
       y_22=> store_value_22,
       y_23=> store_value_23,
       y_24=> store_value_24,
       y_25=> store_value_25,
       y_26=> store_value_26,
       y_27=> store_value_27,
       y_28=> store_value_28,
       y_29=> store_value_29,
       y_30=> store_value_30,
       y_31=> store_value_31,
       y_32=> store_value_32,
       y_33=> store_value_33,
       y_34=> store_value_34,
       y_35=> store_value_35,
       y_36=> store_value_36,
       y_37=> store_value_37,
       y_38=> store_value_38,
       y_39=> store_value_39,
       y_40=> store_value_40,
       y_41=> store_value_41,
       y_42=> store_value_42,
       y_43=> store_value_43,
       y_44=> store_value_44,
       y_45=> store_value_45,
       y_46=> store_value_46,
       y_47=> store_value_47,
       y_48=> store_value_48,
       y_49=> store_value_49,
       y_50=> store_value_50,
       y_51=> store_value_51,
       y_52=> store_value_52,
       y_53=> store_value_53,
       y_54=> store_value_54,
       y_55=> store_value_55,
       y_56=> store_value_56,
       y_57=> store_value_57,
       y_58=> store_value_58,
       y_59=> store_value_59,
       y_60=> store_value_60,
       y_61=> store_value_61,
       y_62=> store_value_62,
       y_63=> store_value_63,
       y_64=> store_value_64,
       y_65=> store_value_65,
       y_66=> store_value_66,
       y_67=> store_value_67,
       y_68=> store_value_68,
       y_69=> store_value_69,
       y_70=> store_value_70,
       y_71=> store_value_71,
       y_72=> store_value_72,
       y_73=> store_value_73,
       y_74=> store_value_74,
       y_75=> store_value_75,
       y_76=> store_value_76,
       y_77=> store_value_77,
       y_78=> store_value_78,
       y_79=> store_value_79,
       y_80=> store_value_80,
       y_81=> store_value_81,
       y_82=> store_value_82,
       y_83=> store_value_83,
       y_84=> store_value_84,
       y_85=> store_value_85,
       y_86=> store_value_86,
       y_87=> store_value_87,
       y_88=> store_value_88,
       y_89=> store_value_89,
       y_90=> store_value_90,
       y_91=> store_value_91,
       y_92=> store_value_92,
       y_93=> store_value_93,
       y_94=> store_value_94,
       y_95=> store_value_95,
       y_96=> store_value_96,
       y_97=> store_value_97,
       y_98=> store_value_98,
       y_99=> store_value_99,
       y_100=> store_value_100,
       y_101=> store_value_101,
       y_102=> store_value_102,
       y_103=> store_value_103,
       y_104=> store_value_104,
       y_105=> store_value_105,
       y_106=> store_value_106,
       y_107=> store_value_107,
       y_108=> store_value_108,
       y_109=> store_value_109,
       y_110=> store_value_110,
       y_111=> store_value_111,
       y_112=> store_value_112,
       y_113=> store_value_113,
       y_114=> store_value_114,
       y_115=> store_value_115,
       y_116=> store_value_116,
       y_117=> store_value_117,
       y_118=> store_value_118,
       y_119=> store_value_119,
       y_120=> store_value_120,
       y_121=> store_value_121,
       y_122=> store_value_122,
       y_123=> store_value_123,
       y_124=> store_value_124,
       y_125=> store_value_125,
       y_126=> store_value_126,
       y_127=> store_value_127,
       y_128=> store_value_128,
       y_129=> store_value_129,
       y_130=> store_value_130,
       y_131=> store_value_131,
       y_132=> store_value_132,
       y_133=> store_value_133,
       y_134=> store_value_134,
       y_135=> store_value_135,
       y_136=> store_value_136,
       y_137=> store_value_137,
       y_138=> store_value_138,
       y_139=> store_value_139,
       y_140=> store_value_140,
       y_141=> store_value_141,
       y_142=> store_value_142,
       y_143=> store_value_143,
       y_144=> store_value_144,
       y_145=> store_value_145,
       y_146=> store_value_146,
       y_147=> store_value_147,
       y_148=> store_value_148,
       y_149=> store_value_149,
       y_150=> store_value_150,
       y_151=> store_value_151,
       y_152=> store_value_152,
       y_153=> store_value_153,
       y_154=> store_value_154,
       y_155=> store_value_155,
       y_156=> store_value_156,
       y_157=> store_value_157,
       y_158=> store_value_158,
       y_159=> store_value_159,
       y_160=> store_value_160,
       y_161=> store_value_161,
       y_162=> store_value_162,
       y_163=> store_value_163,
       y_164=> store_value_164,
       y_165=> store_value_165,
       y_166=> store_value_166,
       y_167=> store_value_167,
       y_168=> store_value_168,
       y_169=> store_value_169,
       y_170=> store_value_170,
       y_171=> store_value_171,
       y_172=> store_value_172,
       y_173=> store_value_173,
       y_174=> store_value_174,
       y_175=> store_value_175,
       y_176=> store_value_176,
       y_177=> store_value_177,
       y_178=> store_value_178,
       y_179=> store_value_179,
       y_180=> store_value_180,
       y_181=> store_value_181,
       y_182=> store_value_182,
       y_183=> store_value_183,
       y_184=> store_value_184,
       y_185=> store_value_185,
       y_186=> store_value_186,
       y_187=> store_value_187,
       y_188=> store_value_188,
       y_189=> store_value_189,
       y_190=> store_value_190,
       y_191=> store_value_191,
       y_192=> store_value_192,
       y_193=> store_value_193,
       y_194=> store_value_194,
       y_195=> store_value_195,
       y_196=> store_value_196,
       y_197=> store_value_197,
       y_198=> store_value_198,
       y_199=> store_value_199,
       y_200=> store_value_200,
       y_201=> store_value_201,
       y_202=> store_value_202,
       y_203=> store_value_203,
       y_204=> store_value_204,
       y_205=> store_value_205,
       y_206=> store_value_206,
       y_207=> store_value_207,
       y_208=> store_value_208,
       y_209=> store_value_209,
       y_210=> store_value_210,
       y_211=> store_value_211,
       y_212=> store_value_212,
       y_213=> store_value_213,
       y_214=> store_value_214,
       y_215=> store_value_215,
       y_216=> store_value_216,
       y_217=> store_value_217,
       y_218=> store_value_218,
       y_219=> store_value_219,
       y_220=> store_value_220,
       y_221=> store_value_221,
       y_222=> store_value_222,
       y_223=> store_value_223,
       y_224=> store_value_224,
       y_225=> store_value_225,
       y_226=> store_value_226,
       y_227=> store_value_227,
       y_228=> store_value_228,
       y_229=> store_value_229,
       y_230=> store_value_230,
       y_231=> store_value_231,
       y_232=> store_value_232,
       y_233=> store_value_233,
       y_234=> store_value_234,
       y_235=> store_value_235,
       y_236=> store_value_236,
       y_237=> store_value_237,
       y_238=> store_value_238,
       y_239=> store_value_239,
       y_240=> store_value_240,
       y_241=> store_value_241,
       y_242=> store_value_242,
       y_243=> store_value_243,
       y_244=> store_value_244,
       y_245=> store_value_245,
       y_246=> store_value_246,
       y_247=> store_value_247,
       y_248=> store_value_248,
       y_249=> store_value_249,
       y_250=> store_value_250,
       y_251=> store_value_251,
       y_252=> store_value_252,
       y_253=> store_value_253,
       y_254=> store_value_254,
       y_255=> store_value_255,
       y_256=> store_value_256,
       y_257=> store_value_257,
       y_258=> store_value_258,
       y_259=> store_value_259,
       y_260=> store_value_260,
       y_261=> store_value_261,
       y_262=> store_value_262,
       y_263=> store_value_263,
       y_264=> store_value_264,
       y_265=> store_value_265,
       y_266=> store_value_266,
       y_267=> store_value_267,
       y_268=> store_value_268,
       y_269=> store_value_269,
       y_270=> store_value_270,
       y_271=> store_value_271,
       y_272=> store_value_272,
       y_273=> store_value_273,
       y_274=> store_value_274,
       y_275=> store_value_275,
       y_276=> store_value_276,
       y_277=> store_value_277,
       y_278=> store_value_278,
       y_279=> store_value_279,
       y_280=> store_value_280,
       y_281=> store_value_281,
       y_282=> store_value_282,
       y_283=> store_value_283,
       y_284=> store_value_284,
       y_285=> store_value_285,
       y_286=> store_value_286,
       y_287=> store_value_287,
       y_288=> store_value_288,
       y_289=> store_value_289,
       y_290=> store_value_290,
       y_291=> store_value_291,
       y_292=> store_value_292,
       y_293=> store_value_293,
       y_294=> store_value_294,
       y_295=> store_value_295,
       y_296=> store_value_296,
       y_297=> store_value_297,
       y_298=> store_value_298,
       y_299=> store_value_299,
       y_300=> store_value_300,
       y_301=> store_value_301,
       y_302=> store_value_302,
       y_303=> store_value_303,
       y_304=> store_value_304,
       y_305=> store_value_305,
       y_306=> store_value_306,
       y_307=> store_value_307,
       y_308=> store_value_308,
       y_309=> store_value_309,
       y_310=> store_value_310,
       y_311=> store_value_311,
       y_312=> store_value_312,
       y_313=> store_value_313,
       y_314=> store_value_314,
       y_315=> store_value_315,
       y_316=> store_value_316,
       y_317=> store_value_317,
       y_318=> store_value_318,
       y_319=> store_value_319,
       y_320=> store_value_320,
       y_321=> store_value_321,
       y_322=> store_value_322,
       y_323=> store_value_323,
       y_324=> store_value_324,
       y_325=> store_value_325,
       y_326=> store_value_326,
       y_327=> store_value_327,
       y_328=> store_value_328,
       y_329=> store_value_329,
       y_330=> store_value_330,
       y_331=> store_value_331,
       y_332=> store_value_332,
       y_333=> store_value_333,
       y_334=> store_value_334,
       y_335=> store_value_335,
       y_336=> store_value_336,
       y_337=> store_value_337,
       y_338=> store_value_338,
       y_339=> store_value_339,
       y_340=> store_value_340,
       y_341=> store_value_341,
       y_342=> store_value_342,
       y_343=> store_value_343,
       y_344=> store_value_344,
       y_345=> store_value_345,
       y_346=> store_value_346,
       y_347=> store_value_347,
       y_348=> store_value_348,
       y_349=> store_value_349,
       y_350=> store_value_350,
       y_351=> store_value_351,
       y_352=> store_value_352,
       y_353=> store_value_353,
       y_354=> store_value_354,
       y_355=> store_value_355,
       y_356=> store_value_356,
       y_357=> store_value_357,
       y_358=> store_value_358,
       y_359=> store_value_359,
       y_360=> store_value_360,
       y_361=> store_value_361,
       y_362=> store_value_362,
       y_363=> store_value_363,
       y_364=> store_value_364,
       y_365=> store_value_365,
       y_366=> store_value_366,
       y_367=> store_value_367,
       y_368=> store_value_368,
       y_369=> store_value_369,
       y_370=> store_value_370,
       y_371=> store_value_371,
       y_372=> store_value_372,
       y_373=> store_value_373,
       y_374=> store_value_374,
       y_375=> store_value_375,
       y_376=> store_value_376,
       y_377=> store_value_377,
       y_378=> store_value_378,
       y_379=> store_value_379,
       y_380=> store_value_380,
       y_381=> store_value_381,
       y_382=> store_value_382,
       y_383=> store_value_383,
       y_384=> store_value_384,
       y_385=> store_value_385,
       y_386=> store_value_386,
       y_387=> store_value_387,
       y_388=> store_value_388,
       y_389=> store_value_389,
       y_390=> store_value_390,
       y_391=> store_value_391,
       y_392=> store_value_392,
       y_393=> store_value_393,
       y_394=> store_value_394,
       y_395=> store_value_395,
       y_396=> store_value_396,
       y_397=> store_value_397,
       y_398=> store_value_398,
       y_399=> store_value_399,
       y_400=> store_value_400,
       y_401=> store_value_401,
       y_402=> store_value_402,
       y_403=> store_value_403,
       y_404=> store_value_404,
       y_405=> store_value_405,
       y_406=> store_value_406,
       y_407=> store_value_407,
       y_408=> store_value_408,
       y_409=> store_value_409,
       y_410=> store_value_410,
       y_411=> store_value_411,
       y_412=> store_value_412,
       y_413=> store_value_413,
       y_414=> store_value_414,
       y_415=> store_value_415,
       y_416=> store_value_416,
       y_417=> store_value_417,
       y_418=> store_value_418,
       y_419=> store_value_419,
       y_420=> store_value_420,
       y_421=> store_value_421,
       y_422=> store_value_422,
       y_423=> store_value_423,
       y_424=> store_value_424,
       y_425=> store_value_425,
       y_426=> store_value_426,
       y_427=> store_value_427,
       y_428=> store_value_428,
       y_429=> store_value_429,
       y_430=> store_value_430,
       y_431=> store_value_431,
       y_432=> store_value_432,
       y_433=> store_value_433,
       y_434=> store_value_434,
       y_435=> store_value_435,
       y_436=> store_value_436,
       y_437=> store_value_437,
       y_438=> store_value_438,
       y_439=> store_value_439,
       y_440=> store_value_440,
       y_441=> store_value_441,
       y_442=> store_value_442,
       y_443=> store_value_443,
       y_444=> store_value_444,
       y_445=> store_value_445,
       y_446=> store_value_446,
       y_447=> store_value_447,
       y_448=> store_value_448,
       y_449=> store_value_449,
       y_450=> store_value_450,
       y_451=> store_value_451,
       y_452=> store_value_452,
       y_453=> store_value_453,
       y_454=> store_value_454,
       y_455=> store_value_455,
       y_456=> store_value_456,
       y_457=> store_value_457,
       y_458=> store_value_458,
       y_459=> store_value_459,
       y_460=> store_value_460,
       y_461=> store_value_461,
       y_462=> store_value_462,
       y_463=> store_value_463,
       y_464=> store_value_464,
       y_465=> store_value_465,
       y_466=> store_value_466,
       y_467=> store_value_467,
       y_468=> store_value_468,
       y_469=> store_value_469,
       y_470=> store_value_470,
       y_471=> store_value_471,
       y_472=> store_value_472,
       y_473=> store_value_473,
       y_474=> store_value_474,
       y_475=> store_value_475,
       y_476=> store_value_476,
       y_477=> store_value_477,
       y_478=> store_value_478,
       y_479=> store_value_479,
       y_480=> store_value_480,
       y_481=> store_value_481,
       y_482=> store_value_482,
       y_483=> store_value_483,
       y_484=> store_value_484,
       y_485=> store_value_485,
       y_486=> store_value_486,
       y_487=> store_value_487,
       y_488=> store_value_488,
       y_489=> store_value_489,
       y_490=> store_value_490,
       y_491=> store_value_491,
       y_492=> store_value_492,
       y_493=> store_value_493,
       y_494=> store_value_494,
       y_495=> store_value_495,
       y_496=> store_value_496,
       y_497=> store_value_497,
       y_498=> store_value_498,
       y_499=> store_value_499,
       y_500=> store_value_500,
       y_501=> store_value_501,
       y_502=> store_value_502,
       y_503=> store_value_503,
       y_504=> store_value_504,
       y_505=> store_value_505,
       y_506=> store_value_506,
       y_507=> store_value_507,
       y_508=> store_value_508,
       y_509=> store_value_509,
       y_510=> store_value_510,
       y_511=> store_value_511,
       y_512=> store_value_512,
       y_513=> store_value_513,
       y_514=> store_value_514,
       y_515=> store_value_515,
       y_516=> store_value_516,
       y_517=> store_value_517,
       y_518=> store_value_518,
       y_519=> store_value_519,
       y_520=> store_value_520,
       y_521=> store_value_521,
       y_522=> store_value_522,
       y_523=> store_value_523,
       y_524=> store_value_524,
       y_525=> store_value_525,
       y_526=> store_value_526,
       y_527=> store_value_527,
       y_528=> store_value_528,
       y_529=> store_value_529,
       y_530=> store_value_530,
       y_531=> store_value_531,
       y_532=> store_value_532,
       y_533=> store_value_533,
       y_534=> store_value_534,
       y_535=> store_value_535,
       y_536=> store_value_536,
       y_537=> store_value_537,
       y_538=> store_value_538,
       y_539=> store_value_539,
       y_540=> store_value_540,
       y_541=> store_value_541,
       y_542=> store_value_542,
       y_543=> store_value_543,
       y_544=> store_value_544,
       y_545=> store_value_545,
       y_546=> store_value_546,
       y_547=> store_value_547,
       y_548=> store_value_548,
       y_549=> store_value_549,
       y_550=> store_value_550,
       y_551=> store_value_551,
       y_552=> store_value_552,
       y_553=> store_value_553,
       y_554=> store_value_554,
       y_555=> store_value_555,
       y_556=> store_value_556,
       y_557=> store_value_557,
       y_558=> store_value_558,
       y_559=> store_value_559,
       y_560=> store_value_560,
       y_561=> store_value_561,
       y_562=> store_value_562,
       y_563=> store_value_563,
       y_564=> store_value_564,
       y_565=> store_value_565,
       y_566=> store_value_566,
       y_567=> store_value_567,
       y_568=> store_value_568,
       y_569=> store_value_569,
       y_570=> store_value_570,
       y_571=> store_value_571,
       y_572=> store_value_572,
       y_573=> store_value_573,
       y_574=> store_value_574,
       y_575=> store_value_575,
       y_576=> store_value_576,
       y_577=> store_value_577,
       y_578=> store_value_578,
       y_579=> store_value_579,
       y_580=> store_value_580,
       y_581=> store_value_581,
       y_582=> store_value_582,
       y_583=> store_value_583,
       y_584=> store_value_584,
       y_585=> store_value_585,
       y_586=> store_value_586,
       y_587=> store_value_587,
       y_588=> store_value_588,
       y_589=> store_value_589,
       y_590=> store_value_590,
       y_591=> store_value_591,
       y_592=> store_value_592,
       y_593=> store_value_593,
       y_594=> store_value_594,
       y_595=> store_value_595,
       y_596=> store_value_596,
       y_597=> store_value_597,
       y_598=> store_value_598,
       y_599=> store_value_599,
       y_600=> store_value_600,
       y_601=> store_value_601,
       y_602=> store_value_602,
       y_603=> store_value_603,
       y_604=> store_value_604,
       y_605=> store_value_605,
       y_606=> store_value_606,
       y_607=> store_value_607,
       y_608=> store_value_608,
       y_609=> store_value_609,
       y_610=> store_value_610,
       y_611=> store_value_611,
       y_612=> store_value_612,
       y_613=> store_value_613,
       y_614=> store_value_614,
       y_615=> store_value_615,
       y_616=> store_value_616,
       y_617=> store_value_617,
       y_618=> store_value_618,
       y_619=> store_value_619,
       y_620=> store_value_620,
       y_621=> store_value_621,
       y_622=> store_value_622,
       y_623=> store_value_623,
       y_624=> store_value_624,
       y_625=> store_value_625,
       y_626=> store_value_626,
       y_627=> store_value_627,
       y_628=> store_value_628,
       y_629=> store_value_629,
       y_630=> store_value_630,
       y_631=> store_value_631,
       y_632=> store_value_632,
       y_633=> store_value_633,
       y_634=> store_value_634,
       y_635=> store_value_635,
       y_636=> store_value_636,
       y_637=> store_value_637,
       y_638=> store_value_638,
       y_639=> store_value_639,
       y_640=> store_value_640,
       y_641=> store_value_641,
       y_642=> store_value_642,
       y_643=> store_value_643,
       y_644=> store_value_644,
       y_645=> store_value_645,
       y_646=> store_value_646,
       y_647=> store_value_647,
       y_648=> store_value_648,
       y_649=> store_value_649,
       y_650=> store_value_650,
       y_651=> store_value_651,
       y_652=> store_value_652,
       y_653=> store_value_653,
       y_654=> store_value_654,
       y_655=> store_value_655,
       y_656=> store_value_656,
       y_657=> store_value_657,
       y_658=> store_value_658,
       y_659=> store_value_659,
       y_660=> store_value_660,
       y_661=> store_value_661,
       y_662=> store_value_662,
       y_663=> store_value_663,
       y_664=> store_value_664,
       y_665=> store_value_665,
       y_666=> store_value_666,
       y_667=> store_value_667,
       y_668=> store_value_668,
       y_669=> store_value_669,
       y_670=> store_value_670,
       y_671=> store_value_671,
       y_672=> store_value_672,
       y_673=> store_value_673,
       y_674=> store_value_674,
       y_675=> store_value_675,
       y_676=> store_value_676,
       y_677=> store_value_677,
       y_678=> store_value_678,
       y_679=> store_value_679,
       y_680=> store_value_680,
       y_681=> store_value_681,
       y_682=> store_value_682,
       y_683=> store_value_683,
       y_684=> store_value_684,
       y_685=> store_value_685,
       y_686=> store_value_686,
       y_687=> store_value_687,
       y_688=> store_value_688,
       y_689=> store_value_689,
       y_690=> store_value_690,
       y_691=> store_value_691,
       y_692=> store_value_692,
       y_693=> store_value_693,
       y_694=> store_value_694,
       y_695=> store_value_695,
       y_696=> store_value_696,
       y_697=> store_value_697,
       y_698=> store_value_698,
       y_699=> store_value_699,
       y_700=> store_value_700,
       y_701=> store_value_701,
       y_702=> store_value_702,
       y_703=> store_value_703,
       y_704=> store_value_704,
       y_705=> store_value_705,
       y_706=> store_value_706,
       y_707=> store_value_707,
       y_708=> store_value_708,
       y_709=> store_value_709,
       y_710=> store_value_710,
       y_711=> store_value_711,
       y_712=> store_value_712,
       y_713=> store_value_713,
       y_714=> store_value_714,
       y_715=> store_value_715,
       y_716=> store_value_716,
       y_717=> store_value_717,
       y_718=> store_value_718,
       y_719=> store_value_719,
       y_720=> store_value_720,
       y_721=> store_value_721,
       y_722=> store_value_722,
       y_723=> store_value_723,
       y_724=> store_value_724,
       y_725=> store_value_725,
       y_726=> store_value_726,
       y_727=> store_value_727,
       y_728=> store_value_728,
       y_729=> store_value_729,
       y_730=> store_value_730,
       y_731=> store_value_731,
       y_732=> store_value_732,
       y_733=> store_value_733,
       y_734=> store_value_734,
       y_735=> store_value_735,
       y_736=> store_value_736,
       y_737=> store_value_737,
       y_738=> store_value_738,
       y_739=> store_value_739,
       y_740=> store_value_740,
       y_741=> store_value_741,
       y_742=> store_value_742,
       y_743=> store_value_743,
       y_744=> store_value_744,
       y_745=> store_value_745,
       y_746=> store_value_746,
       y_747=> store_value_747,
       y_748=> store_value_748,
       y_749=> store_value_749,
       y_750=> store_value_750,
       y_751=> store_value_751,
       y_752=> store_value_752,
       y_753=> store_value_753,
       y_754=> store_value_754,
       y_755=> store_value_755,
       y_756=> store_value_756,
       y_757=> store_value_757,
       y_758=> store_value_758,
       y_759=> store_value_759,
       y_760=> store_value_760,
       y_761=> store_value_761,
       y_762=> store_value_762,
       y_763=> store_value_763,
       y_764=> store_value_764,
       y_765=> store_value_765,
       y_766=> store_value_766,
       y_767=> store_value_767,
       y_768=> store_value_768,
       y_769=> store_value_769,
       y_770=> store_value_770,
       y_771=> store_value_771,
       y_772=> store_value_772,
       y_773=> store_value_773,
       y_774=> store_value_774,
       y_775=> store_value_775,
       y_776=> store_value_776,
       y_777=> store_value_777,
       y_778=> store_value_778,
       y_779=> store_value_779,
       y_780=> store_value_780,
       y_781=> store_value_781,
       y_782=> store_value_782,
       y_783=> store_value_783
		);
   ut0_fully_connected_layer: fully_connected_layer port map(
       clk=> clk,
       x_0=> store_value_0,
       x_1=> store_value_1,
       x_2=> store_value_2,
       x_3=> store_value_3,
       x_4=> store_value_4,
       x_5=> store_value_5,
       x_6=> store_value_6,
       x_7=> store_value_7,
       x_8=> store_value_8,
       x_9=> store_value_9,
       x_10=> store_value_10,
       x_11=> store_value_11,
       x_12=> store_value_12,
       x_13=> store_value_13,
       x_14=> store_value_14,
       x_15=> store_value_15,
       x_16=> store_value_16,
       x_17=> store_value_17,
       x_18=> store_value_18,
       x_19=> store_value_19,
       x_20=> store_value_20,
       x_21=> store_value_21,
       x_22=> store_value_22,
       x_23=> store_value_23,
       x_24=> store_value_24,
       x_25=> store_value_25,
       x_26=> store_value_26,
       x_27=> store_value_27,
       x_28=> store_value_28,
       x_29=> store_value_29,
       x_30=> store_value_30,
       x_31=> store_value_31,
       x_32=> store_value_32,
       x_33=> store_value_33,
       x_34=> store_value_34,
       x_35=> store_value_35,
       x_36=> store_value_36,
       x_37=> store_value_37,
       x_38=> store_value_38,
       x_39=> store_value_39,
       x_40=> store_value_40,
       x_41=> store_value_41,
       x_42=> store_value_42,
       x_43=> store_value_43,
       x_44=> store_value_44,
       x_45=> store_value_45,
       x_46=> store_value_46,
       x_47=> store_value_47,
       x_48=> store_value_48,
       x_49=> store_value_49,
       x_50=> store_value_50,
       x_51=> store_value_51,
       x_52=> store_value_52,
       x_53=> store_value_53,
       x_54=> store_value_54,
       x_55=> store_value_55,
       x_56=> store_value_56,
       x_57=> store_value_57,
       x_58=> store_value_58,
       x_59=> store_value_59,
       x_60=> store_value_60,
       x_61=> store_value_61,
       x_62=> store_value_62,
       x_63=> store_value_63,
       x_64=> store_value_64,
       x_65=> store_value_65,
       x_66=> store_value_66,
       x_67=> store_value_67,
       x_68=> store_value_68,
       x_69=> store_value_69,
       x_70=> store_value_70,
       x_71=> store_value_71,
       x_72=> store_value_72,
       x_73=> store_value_73,
       x_74=> store_value_74,
       x_75=> store_value_75,
       x_76=> store_value_76,
       x_77=> store_value_77,
       x_78=> store_value_78,
       x_79=> store_value_79,
       x_80=> store_value_80,
       x_81=> store_value_81,
       x_82=> store_value_82,
       x_83=> store_value_83,
       x_84=> store_value_84,
       x_85=> store_value_85,
       x_86=> store_value_86,
       x_87=> store_value_87,
       x_88=> store_value_88,
       x_89=> store_value_89,
       x_90=> store_value_90,
       x_91=> store_value_91,
       x_92=> store_value_92,
       x_93=> store_value_93,
       x_94=> store_value_94,
       x_95=> store_value_95,
       x_96=> store_value_96,
       x_97=> store_value_97,
       x_98=> store_value_98,
       x_99=> store_value_99,
       x_100=> store_value_100,
       x_101=> store_value_101,
       x_102=> store_value_102,
       x_103=> store_value_103,
       x_104=> store_value_104,
       x_105=> store_value_105,
       x_106=> store_value_106,
       x_107=> store_value_107,
       x_108=> store_value_108,
       x_109=> store_value_109,
       x_110=> store_value_110,
       x_111=> store_value_111,
       x_112=> store_value_112,
       x_113=> store_value_113,
       x_114=> store_value_114,
       x_115=> store_value_115,
       x_116=> store_value_116,
       x_117=> store_value_117,
       x_118=> store_value_118,
       x_119=> store_value_119,
       x_120=> store_value_120,
       x_121=> store_value_121,
       x_122=> store_value_122,
       x_123=> store_value_123,
       x_124=> store_value_124,
       x_125=> store_value_125,
       x_126=> store_value_126,
       x_127=> store_value_127,
       x_128=> store_value_128,
       x_129=> store_value_129,
       x_130=> store_value_130,
       x_131=> store_value_131,
       x_132=> store_value_132,
       x_133=> store_value_133,
       x_134=> store_value_134,
       x_135=> store_value_135,
       x_136=> store_value_136,
       x_137=> store_value_137,
       x_138=> store_value_138,
       x_139=> store_value_139,
       x_140=> store_value_140,
       x_141=> store_value_141,
       x_142=> store_value_142,
       x_143=> store_value_143,
       x_144=> store_value_144,
       x_145=> store_value_145,
       x_146=> store_value_146,
       x_147=> store_value_147,
       x_148=> store_value_148,
       x_149=> store_value_149,
       x_150=> store_value_150,
       x_151=> store_value_151,
       x_152=> store_value_152,
       x_153=> store_value_153,
       x_154=> store_value_154,
       x_155=> store_value_155,
       x_156=> store_value_156,
       x_157=> store_value_157,
       x_158=> store_value_158,
       x_159=> store_value_159,
       x_160=> store_value_160,
       x_161=> store_value_161,
       x_162=> store_value_162,
       x_163=> store_value_163,
       x_164=> store_value_164,
       x_165=> store_value_165,
       x_166=> store_value_166,
       x_167=> store_value_167,
       x_168=> store_value_168,
       x_169=> store_value_169,
       x_170=> store_value_170,
       x_171=> store_value_171,
       x_172=> store_value_172,
       x_173=> store_value_173,
       x_174=> store_value_174,
       x_175=> store_value_175,
       x_176=> store_value_176,
       x_177=> store_value_177,
       x_178=> store_value_178,
       x_179=> store_value_179,
       x_180=> store_value_180,
       x_181=> store_value_181,
       x_182=> store_value_182,
       x_183=> store_value_183,
       x_184=> store_value_184,
       x_185=> store_value_185,
       x_186=> store_value_186,
       x_187=> store_value_187,
       x_188=> store_value_188,
       x_189=> store_value_189,
       x_190=> store_value_190,
       x_191=> store_value_191,
       x_192=> store_value_192,
       x_193=> store_value_193,
       x_194=> store_value_194,
       x_195=> store_value_195,
       x_196=> store_value_196,
       x_197=> store_value_197,
       x_198=> store_value_198,
       x_199=> store_value_199,
       x_200=> store_value_200,
       x_201=> store_value_201,
       x_202=> store_value_202,
       x_203=> store_value_203,
       x_204=> store_value_204,
       x_205=> store_value_205,
       x_206=> store_value_206,
       x_207=> store_value_207,
       x_208=> store_value_208,
       x_209=> store_value_209,
       x_210=> store_value_210,
       x_211=> store_value_211,
       x_212=> store_value_212,
       x_213=> store_value_213,
       x_214=> store_value_214,
       x_215=> store_value_215,
       x_216=> store_value_216,
       x_217=> store_value_217,
       x_218=> store_value_218,
       x_219=> store_value_219,
       x_220=> store_value_220,
       x_221=> store_value_221,
       x_222=> store_value_222,
       x_223=> store_value_223,
       x_224=> store_value_224,
       x_225=> store_value_225,
       x_226=> store_value_226,
       x_227=> store_value_227,
       x_228=> store_value_228,
       x_229=> store_value_229,
       x_230=> store_value_230,
       x_231=> store_value_231,
       x_232=> store_value_232,
       x_233=> store_value_233,
       x_234=> store_value_234,
       x_235=> store_value_235,
       x_236=> store_value_236,
       x_237=> store_value_237,
       x_238=> store_value_238,
       x_239=> store_value_239,
       x_240=> store_value_240,
       x_241=> store_value_241,
       x_242=> store_value_242,
       x_243=> store_value_243,
       x_244=> store_value_244,
       x_245=> store_value_245,
       x_246=> store_value_246,
       x_247=> store_value_247,
       x_248=> store_value_248,
       x_249=> store_value_249,
       x_250=> store_value_250,
       x_251=> store_value_251,
       x_252=> store_value_252,
       x_253=> store_value_253,
       x_254=> store_value_254,
       x_255=> store_value_255,
       x_256=> store_value_256,
       x_257=> store_value_257,
       x_258=> store_value_258,
       x_259=> store_value_259,
       x_260=> store_value_260,
       x_261=> store_value_261,
       x_262=> store_value_262,
       x_263=> store_value_263,
       x_264=> store_value_264,
       x_265=> store_value_265,
       x_266=> store_value_266,
       x_267=> store_value_267,
       x_268=> store_value_268,
       x_269=> store_value_269,
       x_270=> store_value_270,
       x_271=> store_value_271,
       x_272=> store_value_272,
       x_273=> store_value_273,
       x_274=> store_value_274,
       x_275=> store_value_275,
       x_276=> store_value_276,
       x_277=> store_value_277,
       x_278=> store_value_278,
       x_279=> store_value_279,
       x_280=> store_value_280,
       x_281=> store_value_281,
       x_282=> store_value_282,
       x_283=> store_value_283,
       x_284=> store_value_284,
       x_285=> store_value_285,
       x_286=> store_value_286,
       x_287=> store_value_287,
       x_288=> store_value_288,
       x_289=> store_value_289,
       x_290=> store_value_290,
       x_291=> store_value_291,
       x_292=> store_value_292,
       x_293=> store_value_293,
       x_294=> store_value_294,
       x_295=> store_value_295,
       x_296=> store_value_296,
       x_297=> store_value_297,
       x_298=> store_value_298,
       x_299=> store_value_299,
       x_300=> store_value_300,
       x_301=> store_value_301,
       x_302=> store_value_302,
       x_303=> store_value_303,
       x_304=> store_value_304,
       x_305=> store_value_305,
       x_306=> store_value_306,
       x_307=> store_value_307,
       x_308=> store_value_308,
       x_309=> store_value_309,
       x_310=> store_value_310,
       x_311=> store_value_311,
       x_312=> store_value_312,
       x_313=> store_value_313,
       x_314=> store_value_314,
       x_315=> store_value_315,
       x_316=> store_value_316,
       x_317=> store_value_317,
       x_318=> store_value_318,
       x_319=> store_value_319,
       x_320=> store_value_320,
       x_321=> store_value_321,
       x_322=> store_value_322,
       x_323=> store_value_323,
       x_324=> store_value_324,
       x_325=> store_value_325,
       x_326=> store_value_326,
       x_327=> store_value_327,
       x_328=> store_value_328,
       x_329=> store_value_329,
       x_330=> store_value_330,
       x_331=> store_value_331,
       x_332=> store_value_332,
       x_333=> store_value_333,
       x_334=> store_value_334,
       x_335=> store_value_335,
       x_336=> store_value_336,
       x_337=> store_value_337,
       x_338=> store_value_338,
       x_339=> store_value_339,
       x_340=> store_value_340,
       x_341=> store_value_341,
       x_342=> store_value_342,
       x_343=> store_value_343,
       x_344=> store_value_344,
       x_345=> store_value_345,
       x_346=> store_value_346,
       x_347=> store_value_347,
       x_348=> store_value_348,
       x_349=> store_value_349,
       x_350=> store_value_350,
       x_351=> store_value_351,
       x_352=> store_value_352,
       x_353=> store_value_353,
       x_354=> store_value_354,
       x_355=> store_value_355,
       x_356=> store_value_356,
       x_357=> store_value_357,
       x_358=> store_value_358,
       x_359=> store_value_359,
       x_360=> store_value_360,
       x_361=> store_value_361,
       x_362=> store_value_362,
       x_363=> store_value_363,
       x_364=> store_value_364,
       x_365=> store_value_365,
       x_366=> store_value_366,
       x_367=> store_value_367,
       x_368=> store_value_368,
       x_369=> store_value_369,
       x_370=> store_value_370,
       x_371=> store_value_371,
       x_372=> store_value_372,
       x_373=> store_value_373,
       x_374=> store_value_374,
       x_375=> store_value_375,
       x_376=> store_value_376,
       x_377=> store_value_377,
       x_378=> store_value_378,
       x_379=> store_value_379,
       x_380=> store_value_380,
       x_381=> store_value_381,
       x_382=> store_value_382,
       x_383=> store_value_383,
       x_384=> store_value_384,
       x_385=> store_value_385,
       x_386=> store_value_386,
       x_387=> store_value_387,
       x_388=> store_value_388,
       x_389=> store_value_389,
       x_390=> store_value_390,
       x_391=> store_value_391,
       x_392=> store_value_392,
       x_393=> store_value_393,
       x_394=> store_value_394,
       x_395=> store_value_395,
       x_396=> store_value_396,
       x_397=> store_value_397,
       x_398=> store_value_398,
       x_399=> store_value_399,
       x_400=> store_value_400,
       x_401=> store_value_401,
       x_402=> store_value_402,
       x_403=> store_value_403,
       x_404=> store_value_404,
       x_405=> store_value_405,
       x_406=> store_value_406,
       x_407=> store_value_407,
       x_408=> store_value_408,
       x_409=> store_value_409,
       x_410=> store_value_410,
       x_411=> store_value_411,
       x_412=> store_value_412,
       x_413=> store_value_413,
       x_414=> store_value_414,
       x_415=> store_value_415,
       x_416=> store_value_416,
       x_417=> store_value_417,
       x_418=> store_value_418,
       x_419=> store_value_419,
       x_420=> store_value_420,
       x_421=> store_value_421,
       x_422=> store_value_422,
       x_423=> store_value_423,
       x_424=> store_value_424,
       x_425=> store_value_425,
       x_426=> store_value_426,
       x_427=> store_value_427,
       x_428=> store_value_428,
       x_429=> store_value_429,
       x_430=> store_value_430,
       x_431=> store_value_431,
       x_432=> store_value_432,
       x_433=> store_value_433,
       x_434=> store_value_434,
       x_435=> store_value_435,
       x_436=> store_value_436,
       x_437=> store_value_437,
       x_438=> store_value_438,
       x_439=> store_value_439,
       x_440=> store_value_440,
       x_441=> store_value_441,
       x_442=> store_value_442,
       x_443=> store_value_443,
       x_444=> store_value_444,
       x_445=> store_value_445,
       x_446=> store_value_446,
       x_447=> store_value_447,
       x_448=> store_value_448,
       x_449=> store_value_449,
       x_450=> store_value_450,
       x_451=> store_value_451,
       x_452=> store_value_452,
       x_453=> store_value_453,
       x_454=> store_value_454,
       x_455=> store_value_455,
       x_456=> store_value_456,
       x_457=> store_value_457,
       x_458=> store_value_458,
       x_459=> store_value_459,
       x_460=> store_value_460,
       x_461=> store_value_461,
       x_462=> store_value_462,
       x_463=> store_value_463,
       x_464=> store_value_464,
       x_465=> store_value_465,
       x_466=> store_value_466,
       x_467=> store_value_467,
       x_468=> store_value_468,
       x_469=> store_value_469,
       x_470=> store_value_470,
       x_471=> store_value_471,
       x_472=> store_value_472,
       x_473=> store_value_473,
       x_474=> store_value_474,
       x_475=> store_value_475,
       x_476=> store_value_476,
       x_477=> store_value_477,
       x_478=> store_value_478,
       x_479=> store_value_479,
       x_480=> store_value_480,
       x_481=> store_value_481,
       x_482=> store_value_482,
       x_483=> store_value_483,
       x_484=> store_value_484,
       x_485=> store_value_485,
       x_486=> store_value_486,
       x_487=> store_value_487,
       x_488=> store_value_488,
       x_489=> store_value_489,
       x_490=> store_value_490,
       x_491=> store_value_491,
       x_492=> store_value_492,
       x_493=> store_value_493,
       x_494=> store_value_494,
       x_495=> store_value_495,
       x_496=> store_value_496,
       x_497=> store_value_497,
       x_498=> store_value_498,
       x_499=> store_value_499,
       x_500=> store_value_500,
       x_501=> store_value_501,
       x_502=> store_value_502,
       x_503=> store_value_503,
       x_504=> store_value_504,
       x_505=> store_value_505,
       x_506=> store_value_506,
       x_507=> store_value_507,
       x_508=> store_value_508,
       x_509=> store_value_509,
       x_510=> store_value_510,
       x_511=> store_value_511,
       x_512=> store_value_512,
       x_513=> store_value_513,
       x_514=> store_value_514,
       x_515=> store_value_515,
       x_516=> store_value_516,
       x_517=> store_value_517,
       x_518=> store_value_518,
       x_519=> store_value_519,
       x_520=> store_value_520,
       x_521=> store_value_521,
       x_522=> store_value_522,
       x_523=> store_value_523,
       x_524=> store_value_524,
       x_525=> store_value_525,
       x_526=> store_value_526,
       x_527=> store_value_527,
       x_528=> store_value_528,
       x_529=> store_value_529,
       x_530=> store_value_530,
       x_531=> store_value_531,
       x_532=> store_value_532,
       x_533=> store_value_533,
       x_534=> store_value_534,
       x_535=> store_value_535,
       x_536=> store_value_536,
       x_537=> store_value_537,
       x_538=> store_value_538,
       x_539=> store_value_539,
       x_540=> store_value_540,
       x_541=> store_value_541,
       x_542=> store_value_542,
       x_543=> store_value_543,
       x_544=> store_value_544,
       x_545=> store_value_545,
       x_546=> store_value_546,
       x_547=> store_value_547,
       x_548=> store_value_548,
       x_549=> store_value_549,
       x_550=> store_value_550,
       x_551=> store_value_551,
       x_552=> store_value_552,
       x_553=> store_value_553,
       x_554=> store_value_554,
       x_555=> store_value_555,
       x_556=> store_value_556,
       x_557=> store_value_557,
       x_558=> store_value_558,
       x_559=> store_value_559,
       x_560=> store_value_560,
       x_561=> store_value_561,
       x_562=> store_value_562,
       x_563=> store_value_563,
       x_564=> store_value_564,
       x_565=> store_value_565,
       x_566=> store_value_566,
       x_567=> store_value_567,
       x_568=> store_value_568,
       x_569=> store_value_569,
       x_570=> store_value_570,
       x_571=> store_value_571,
       x_572=> store_value_572,
       x_573=> store_value_573,
       x_574=> store_value_574,
       x_575=> store_value_575,
       x_576=> store_value_576,
       x_577=> store_value_577,
       x_578=> store_value_578,
       x_579=> store_value_579,
       x_580=> store_value_580,
       x_581=> store_value_581,
       x_582=> store_value_582,
       x_583=> store_value_583,
       x_584=> store_value_584,
       x_585=> store_value_585,
       x_586=> store_value_586,
       x_587=> store_value_587,
       x_588=> store_value_588,
       x_589=> store_value_589,
       x_590=> store_value_590,
       x_591=> store_value_591,
       x_592=> store_value_592,
       x_593=> store_value_593,
       x_594=> store_value_594,
       x_595=> store_value_595,
       x_596=> store_value_596,
       x_597=> store_value_597,
       x_598=> store_value_598,
       x_599=> store_value_599,
       x_600=> store_value_600,
       x_601=> store_value_601,
       x_602=> store_value_602,
       x_603=> store_value_603,
       x_604=> store_value_604,
       x_605=> store_value_605,
       x_606=> store_value_606,
       x_607=> store_value_607,
       x_608=> store_value_608,
       x_609=> store_value_609,
       x_610=> store_value_610,
       x_611=> store_value_611,
       x_612=> store_value_612,
       x_613=> store_value_613,
       x_614=> store_value_614,
       x_615=> store_value_615,
       x_616=> store_value_616,
       x_617=> store_value_617,
       x_618=> store_value_618,
       x_619=> store_value_619,
       x_620=> store_value_620,
       x_621=> store_value_621,
       x_622=> store_value_622,
       x_623=> store_value_623,
       x_624=> store_value_624,
       x_625=> store_value_625,
       x_626=> store_value_626,
       x_627=> store_value_627,
       x_628=> store_value_628,
       x_629=> store_value_629,
       x_630=> store_value_630,
       x_631=> store_value_631,
       x_632=> store_value_632,
       x_633=> store_value_633,
       x_634=> store_value_634,
       x_635=> store_value_635,
       x_636=> store_value_636,
       x_637=> store_value_637,
       x_638=> store_value_638,
       x_639=> store_value_639,
       x_640=> store_value_640,
       x_641=> store_value_641,
       x_642=> store_value_642,
       x_643=> store_value_643,
       x_644=> store_value_644,
       x_645=> store_value_645,
       x_646=> store_value_646,
       x_647=> store_value_647,
       x_648=> store_value_648,
       x_649=> store_value_649,
       x_650=> store_value_650,
       x_651=> store_value_651,
       x_652=> store_value_652,
       x_653=> store_value_653,
       x_654=> store_value_654,
       x_655=> store_value_655,
       x_656=> store_value_656,
       x_657=> store_value_657,
       x_658=> store_value_658,
       x_659=> store_value_659,
       x_660=> store_value_660,
       x_661=> store_value_661,
       x_662=> store_value_662,
       x_663=> store_value_663,
       x_664=> store_value_664,
       x_665=> store_value_665,
       x_666=> store_value_666,
       x_667=> store_value_667,
       x_668=> store_value_668,
       x_669=> store_value_669,
       x_670=> store_value_670,
       x_671=> store_value_671,
       x_672=> store_value_672,
       x_673=> store_value_673,
       x_674=> store_value_674,
       x_675=> store_value_675,
       x_676=> store_value_676,
       x_677=> store_value_677,
       x_678=> store_value_678,
       x_679=> store_value_679,
       x_680=> store_value_680,
       x_681=> store_value_681,
       x_682=> store_value_682,
       x_683=> store_value_683,
       x_684=> store_value_684,
       x_685=> store_value_685,
       x_686=> store_value_686,
       x_687=> store_value_687,
       x_688=> store_value_688,
       x_689=> store_value_689,
       x_690=> store_value_690,
       x_691=> store_value_691,
       x_692=> store_value_692,
       x_693=> store_value_693,
       x_694=> store_value_694,
       x_695=> store_value_695,
       x_696=> store_value_696,
       x_697=> store_value_697,
       x_698=> store_value_698,
       x_699=> store_value_699,
       x_700=> store_value_700,
       x_701=> store_value_701,
       x_702=> store_value_702,
       x_703=> store_value_703,
       x_704=> store_value_704,
       x_705=> store_value_705,
       x_706=> store_value_706,
       x_707=> store_value_707,
       x_708=> store_value_708,
       x_709=> store_value_709,
       x_710=> store_value_710,
       x_711=> store_value_711,
       x_712=> store_value_712,
       x_713=> store_value_713,
       x_714=> store_value_714,
       x_715=> store_value_715,
       x_716=> store_value_716,
       x_717=> store_value_717,
       x_718=> store_value_718,
       x_719=> store_value_719,
       x_720=> store_value_720,
       x_721=> store_value_721,
       x_722=> store_value_722,
       x_723=> store_value_723,
       x_724=> store_value_724,
       x_725=> store_value_725,
       x_726=> store_value_726,
       x_727=> store_value_727,
       x_728=> store_value_728,
       x_729=> store_value_729,
       x_730=> store_value_730,
       x_731=> store_value_731,
       x_732=> store_value_732,
       x_733=> store_value_733,
       x_734=> store_value_734,
       x_735=> store_value_735,
       x_736=> store_value_736,
       x_737=> store_value_737,
       x_738=> store_value_738,
       x_739=> store_value_739,
       x_740=> store_value_740,
       x_741=> store_value_741,
       x_742=> store_value_742,
       x_743=> store_value_743,
       x_744=> store_value_744,
       x_745=> store_value_745,
       x_746=> store_value_746,
       x_747=> store_value_747,
       x_748=> store_value_748,
       x_749=> store_value_749,
       x_750=> store_value_750,
       x_751=> store_value_751,
       x_752=> store_value_752,
       x_753=> store_value_753,
       x_754=> store_value_754,
       x_755=> store_value_755,
       x_756=> store_value_756,
       x_757=> store_value_757,
       x_758=> store_value_758,
       x_759=> store_value_759,
       x_760=> store_value_760,
       x_761=> store_value_761,
       x_762=> store_value_762,
       x_763=> store_value_763,
       x_764=> store_value_764,
       x_765=> store_value_765,
       x_766=> store_value_766,
       x_767=> store_value_767,
       x_768=> store_value_768,
       x_769=> store_value_769,
       x_770=> store_value_770,
       x_771=> store_value_771,
       x_772=> store_value_772,
       x_773=> store_value_773,
       x_774=> store_value_774,
       x_775=> store_value_775,
       x_776=> store_value_776,
       x_777=> store_value_777,
       x_778=> store_value_778,
       x_779=> store_value_779,
       x_780=> store_value_780,
       x_781=> store_value_781,
       x_782=> store_value_782,
       x_783=> store_value_783,
       y => y
		);
end Behavioral;