library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_3 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_3;

architecture syn of ram_3 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"0000000101110001","1000000000000110","0000000110111111","1000000010101100","1000000000101100","1000000011011001","0000000000011101","0000000011100010","1000000001010111","0000000101101110","0000000111111011","1000000001000111","1000010111110110","1000011011110110","1000001011000010","1000000010000110","1000000101010110","1000000011001101","1000000000110111","1000000100000010","1000000111110110","0000000011010111","0000000011111111","1000000011010111","0000000110011010","0000000011000110","1000000001111100","1000000001000101","0000000011100100","0000000010011011","1000000011010001","1000000011100001","0000000001010000","1000000000000010","1000000000110001","1000001100101000","1000001100101011","1000001100101011","1000111100110011","1001000001011000","1001100000111111","1001101011110101","1001000010111001","1001001100010101","1001101010110001","1001011111011010","1001000011001111","1001011011111011","1001000001110101","1000110111110000","1000000101001110","1000000101011111","1000000100000000","0000000000000110","0000000010110100","0000000111110111","0000000111011101","0000000010110000","1000000011110101","1000001000001110","1000010000010001","1000110000100111","1000111101111001","1001011111001000","1001110100000001","1011001111000111","1000011010101111","0000010000001110","0000001110001001","1000001101001011","1000011110101001","1001001011100110","1001000110100110","1001000100011000","1001001000001100","1001111011111111","1010011110010011","1010000001000011","1001100001101100","1001100000110011","1000100101010100","1000000011100101","1000000011101101","0000000010010100","1000000110100010","1000000000001111","1001000101000001","1001000101101011","1000011001001010","0000110100011100","0000100101001100","0000111111100110","0000111001100001","1000010000110001","1000001010110000","0000100011001011","0000111011000001","0000001101001101","0000110000111110","0000110010000110","0000101100010010","0000101001111110","0000011001100001","1000010110110100","0000011000101001","1000010000011010","1001111100001001","1010100111001011","1001001001111111","1000100011011010","1000000101000100","1000000000111001","0000000110011111","0000101100000000","1000010101111110","0000111101111001","0000001010011011","0000100100011010","0000010110101011","0000011110010001","0000100111101001","1000001101010111","0000010011001110","0000010111110111","0000001001110110","0000001110011011","0000000101100101","0000010000100001","0000001000110000","1000010111000100","0000000101001111","1000000011010000","1000111111101101","1000110011000011","1000001110001000","1001110011111010","1011011001101101","1001010000110110","1000001100111001","1000000110001001","1000000000001001","0000000000100110","1000010110010101","0000001100010011","0000101110001111","0000101101000010","0000010001001010","0000010011110011","0000001100110010","0000000110111001","0000001001110010","1000010010111101","1000010101001101","1000011011011011","1000011100010100","0000000110100101","0000000111001110","1000100111001100","1000011111000100","0000000010100011","1000100101000100","1000011111111010","1000011011110010","1000111001010101","1001011000100000","1011010101111011","1001001011011001","1000010101011101","1000000001000001","0000101110001010","0000001110011011","0000010000100110","1000000101001100","0000011110110111","0000010110000111","0000001000110001","0000100011001110","0000001000111011","0000010011000010","1000001001000111","1000011000001010","0000000100011010","1000000100000100","0000001000010000","0000001000011101","1000011110000011","0000000001001000","1000011101000110","1000100010100101","1000000111010100","1000011001011010","1000100011001110","1000110100010000","1100000000000110","1001000001000110","1000010101010000","1000010111010100","0001001110010101","1000011101011011","1000001011101111","0000101001001111","0000100000101100","0000011101000111","1000000011101000","0000001101000011","0000000011001010","1000010110011000","1000100001001111","1000001110101011","1000100011010000","0000001100001000","0000000011000011","1000010001111111","1000010010001001","1000100010010011","1000010000011011","1000000010011010","1000011110101111","1000101100010010","1000000111111001","1000110111100110","1100101010000010","1001001010100000","1000011001010000","1000101001000000","1001100111100110","1000001100111000","1000001101110100","0000001111011100","0000000010110100","0000001000011110","1000011100011000","1000010101001000","1000010111100101","1000010100100001","1000010100001111","1000011011001110","1000100010110001","1000010110000011","1000000000000100","1000001011100001","1000010001011100","0000000111011010","1000001010010110","1000001100100110","1000010000100100","1000000101111100","1000111011010101","1010010011110101","1100011110000000","1001001011000010","1000000101101111","1000101000010101","1000111110000100","0000101111000001","0000011011010011","0001000001011000","0000001100110111","0000011001011100","1000000000000110","0000001001000011","1000001111011111","1000100110011101","1001001100111110","1001001010111101","1000101111001110","0000000000110001","0000011100000110","0000010000101000","0000001110001001","1000001001010100","1000000001011101","0000000110100100","1000000100100000","1000001001101111","1000010111000011","1010100011110010","1000100101001000","1001110100100101","1000011001100010","1000101001000110","1001011001010000","0000001110011001","0000001100111011","0000000001111000","1000001011110111","0000011001100111","1000010010110111","1000011101011010","1001001101010101","1001011111000001","1001100011010111","1001100010111110","1000011010111100","0000000111011011","0000000110111011","0000001000011111","0000001001011101","0000000110110101","0000000101011100","0000000110001011","0000000000111110","1000000001100101","1000001000000101","1011001101000101","0000010011011100","1010011010010110","1000101011110111","1000101111001100","1000101011111001","1000000011100100","0001000110011111","0000100010010111","1000010100010011","1000000000111011","1001010101010111","1001010110101101","1001010110001100","1001011101110001","1000110101100111","1000100010000000","1000010111110100","0000001111110000","0000001001011110","1000010111000101","0000001110000101","0000000100110011","0000000001000010","0000001001000101","1000000100011100","1000110011011001","1000101100000011","1001011111110010","0000001101010100","1001101000101101","1000110110010011","1000011110101110","1000110111100011","1001100010000010","0000001111000110","1000000110111010","1000110101000001","1001001101010000","1000010010010101","1000110110010011","1000100001110010","1000001010100010","1000011111100001","1000001000010001","1000001101011000","0000100011110110","1000001011111011","1000000110001011","1000001000001001","1000000010100110","1000100101011001","1000011111100100","1001010000111010","1010001000110001","1001001011110001","1000110011000100","0001001011101000","1001000100110011","1000110001111110","1000101110111000","1001000101100111","1010100010100101","0000011001001111","0000000000111100","1000001101111011","1000010101010111","1000101011111001","1000001000111011","1000011001100110","1000011110010110","1000100110111101","1000010000100000","0000001001100100","0000000001110000","1000011110100111","1000001010001000","1000000000011001","0000000110100110","1000011001001010","1000110101101110","1000111101111111","1010000001110000","1000011011011000","1001110111010011","0000001000010011","1001010111011010","1000101101101101","1000110000110010","0001001101001100","0000001001110010","0000000111101101","1000001100100011","1001001010010000","1000011001010000","1000110001011100","1000001111010101","1000010101111100","1000110010011110","1000100001110111","1000000101100110","1000010110110101","1000001100110010","1000010010101011","1000010011100110","1000001010010111","1000001000001101","1000001110000000","1000100110001101","0000000100011101","1000111001011010","1000011111101010","1000100000111101","1001000111001111","1001110010000100","1000101110101110","1000110110110101","0000110010110110","0001001011100111","0000001011010010","1000000011101010","1000000111000011","1000001100010100","1000011111000010","1000010000101001","1000101011100001","1000101111110010","1000010101001100","1000000101000001","1000011010100101","1000000101110000","0000000010010110","1000011011010011","1000001100101100","1000010011100100","0000000010010110","0000010111110111","0000000100110100","0000000011011111","0000001110110000","0000000111100110","1001101111001010","0000111001010101","1000101100001111","1000011000110001","0001000111100000","0000010111010111","0000101100001010","0000011000001001","0000100101101101","1000010111100110","1000101110100101","1000100100001101","1000010011111100","1000110101101000","1000011010011010","1000001001010110","1000000100110001","1000011010011100","1000100100100000","1000101110110000","1000011011000100","0000001001010100","0000001011000111","0000000111000011","1000001100011011","0000000011010110","0000000000001011","0001100110010001","1010100110001111","1000000011101101","1000110111111100","1000000000010011","0001000000111111","1000010100101011","0000011100010101","0000100000000111","0000001111011011","0000000001111001","1000000100000100","1000101001110011","1001010001110011","1001101101011010","1001010111000100","1001000001011011","1001001100111111","1001011000111001","1001000001100101","1000010110000110","0000010001001111","1000001111001110","0000100011010100","1000011001101010","1000010010101111","0000011010000100","1000100111001100","1000011000011100","1011001001000000","1010010010100101","1001000010000011","1001010110011011","0000111000100100","0000001111110110","0000111000001001","0000010111110000","0000011000100110","0000001101110001","1000000001111110","1000000011011001","1000101010110000","1001010011001110","1001100111100111","1001100010110010","1001101011110110","1001010011010110","1000001010111011","0000001011000000","0000010111011101","1000000010010011","0000000111001111","1000001111000110","0000000100101010","0000001111000100","0000001010101101","1000110111000110","1100010010111001","1010000110001011","1000111111000000","1000011100100011","1000101100101000","1000001100101100","0000110100000010","0000011010000011","0000100100001101","0000000001111001","0000001011110110","1000001010111000","1000000000010010","1000011100001100","1001001001101000","1001000001101100","1000111010101000","1000011101101101","1000001001011101","1000000011000001","0000011110110010","0000010011010101","0000001011000011","1000001101110100","0000000011010011","1000011000010111","1000011110001111","1000010000111011","1001011010001110","1010110100001100","1000110110011101","1000000110101101","1000101111110010","1000101011010001","0000110000100111","0000011100000011","0000001101100000","0000100000001110","0000011001100001","0000000011010000","0000010111100000","1000010100100010","1000100110101001","1001001000000001","1000100111111100","1000000100010000","1000001101001010","1000000010110110","0000010110101000","0000010111000010","1000000011101000","0000011000011000","1000000111010011","1000000010010111","0000010110101100","1000000010010000","1001000101101001","0000011111111101","1000100010100110","1000100010100001","0000011010111110","0000100111000000","0000010010000110","0000100101000110","0000000111010100","0000011101010001","0000001111111110","0000000000011101","1000001110010010","1000011011001100","1000100000000000","1000101101100110","1000011100100010","1000011001100010","1000001000111010","0000000101001001","0000000111101110","0000011111010001","0000000010100010","0000000001010001","1000111000000101","1001001001001111","0000001110111100","1010001100000101","1010111110101111","0000001101001001","1000001110000101","1000101011101100","1000011011111110","0000001111101101","0000000110100110","0000011000000111","1000001010100111","0000101011101011","0000000100000010","0000000100000000","1000001010101010","1000001100100000","1000000111010111","1000101110001010","1000101011001100","1000011100111111","0000000000000101","0000000001000101","0000001101100010","1000001011011110","0000001101111111","1000000010110001","1000000010110101","1000110001100000","0000000010111111","1010000101110110","1001000010110000","0000010110101010","1000010000100111","1000000110101101","1000000001110101","0000100111001010","0000100010000110","0000100111110010","0000101011100010","0000010100001100","0000010111101001","0000001011011101","0000000111100010","1000000100110111","0000000010010010","1000100001011011","1000001001000011","1000010100010011","1000001001001001","1000011010010111","0000010000101101","0000011010101100","0000000101000001","1000001111000010","1000011110011010","1001110000101001","1000110100010000","1000010010100010","0000011010000000","0000101011000110","1000000011100000","1000000000010100","0000000000101011","0000011010100000","0001100011010110","0000000001101110","0000011111111010","0000101111000000","0000101101110010","0000011100011011","1000010110111000","0000011000001110","0000011010010101","0000010100011100","0000011111100011","0000001101110010","1000000110000010","0000100011001101","0000100110000000","1000011100011011","1001000000110100","1000111010000010","1000110110111100","1000111101010111","1000010100100010","1001000110011100","1001010100111000","1000010000001100","1000000111011000","0000000111111000","0000000001000100","0001000010010111","1001011001100001","0000001101010110","0000000110100011","0000111000001101","0001000010000111","0001000111001001","0000111100101111","0000100011000100","0001000010000011","0001101100111111","0001000101100010","0000010110001010","1000000001010001","0000011111100111","0000010010001110","0000001100110000","0000110010010011","0000010101110111","1000111111100100","1000110110001110","1010111001100101","1001000101010110","1000101001110100","1000000000100111","0000000011110001","1000000011110110","1000000001010101","0000000001101100","1000110001110101","1000100011101110","1000001111001111","1001001010011100","1000010100110111","1000100000111101","1001000111101100","1000001000111001","1000100111011100","1000101110010011","0000000001110101","1000010011010110","1000010111101101","0000011111011100","0000011001100101","1000000111100011","1000000011110000","1000000010100000","1000010110100101","1000101001101010","1001100101000111","1000001000111010","1000001100101011","1000000110110101","0000000001011111","0000000011100101","1000000001110100","1000000010101001","0000000100111100","1000000101101010","1000000110100001","1000110010010001","1000111110111101","1001011101101101","1010001010010110","1010001101101000","1011011100101000","1010000001000001","1010101001100000","1001101111101110","1100010011101000","1011001011001111","1011111110110110","1010001100011011","1001011110001011","1001110001110001","1001000100001010","1001000111110110","1000011010101110","1000000000111001","0000000011010011","0000000111000101","1000000010001000");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
