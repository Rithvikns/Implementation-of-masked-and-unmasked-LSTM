library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_9 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_9;

architecture syn of ram_9 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"1000000100111011","1000000001100011","0000000101001101","0000000010010000","1000000011011101","1000000111001111","1000000001110010","1000000010101000","1000000101010001","1000000010001100","1000000100110111","0000000110101111","1000010001101110","1000011100110110","0000000001101100","1000000110101000","1000000000100001","1000000111011011","1000000010001100","0000000111001010","0000000111100110","1000000110001101","1000000010100000","0000000111101011","0000000010100010","0000000001000100","1000000010000111","1000000000110011","0000000101001110","0000000011011110","1000000110010101","0000000010000100","1000000110100101","0000000000111010","1000001011101010","1000001101011011","1000001111101000","1000001100100010","1000110101010100","1001001111100011","1001001000111010","1001001111100000","1001001010110010","1001000110110111","1001000000011100","1001001010001101","1001011110011001","1001101011110011","1001001100011000","1001001000011001","1000110011010111","1000100011011100","1000000010000111","1000000101001011","1000000000101000","0000000001110100","0000000100011000","1000000011100010","1000000011011000","1000110110000011","1000110101010111","1000001111011110","1000001110100011","1000111010101001","1000110100011101","1001001000110101","1010010001100011","1001110101011000","1010000011110001","1010011000110101","1100111001000111","1100100010101110","1010010010011111","1011011000000000","1011001101101010","1010101100101111","1001111010110110","1001000110000110","1000110111001000","1000110101100111","1000001001011000","1000000101011111","1000000000110001","0000000111111010","1000000111001111","1000000100011101","1000001110110111","1000111110100010","1000110000111101","1000110110101101","1001001000110111","1001011000101100","1001101011000010","1001100100101101","1011111110101111","1100110010000101","1101011110111111","1101111111110011","1101010111101101","1101100101101001","1110000001011011","1011000011001111","1000001000010101","1000001010011001","1001110111111011","1001110010011111","1001110101011111","1000111101001011","1000011000001111","1000001101101111","1000000000110011","1000000001011010","1000000101111100","0000000100100000","1000000000011101","1000101110000100","1000111110100000","1001010111011110","1001100111110111","1010110101111111","1011001001101010","1100000100111101","1011101011110001","1010001011010101","1001111100001001","1001101011101100","1010001011001001","1010000001101100","1010011011000001","1010000101100111","1001100100011010","1011111010111111","1100100100110101","1100011111001100","1011100000011010","1010101010001001","1001001111010010","1000111110001100","1000100011100010","1000010110001110","1000000011010001","0000000010101111","1000001100010010","1000111111110000","1001110010000110","1011101101100110","1011100011011101","1001011000000001","1001011011101101","1001000010011000","1000101101001011","0000001110111011","1000001001110101","1000000011100101","1000010101011001","1000011010001111","1001101110111101","1001001111010010","1000111110100000","1000010110111000","1000101111011100","1001011010101100","1001000100111010","1011101010101101","1101001010110110","1011000110001110","1001010110100110","1000000000100010","0000000001011000","1000101100001010","1001001100010000","1001111001011110","1000010100111100","1001010111110100","1000010110010010","1001010010111011","1000010011100110","1000000111100110","0000000000001100","0000000100110100","0000001001110110","0000100101110100","0000100011011111","0000000000111010","0000101001101101","0000110001111011","0000100010101011","1000001010010111","1000001100001110","1000011010010001","1000100000000101","1000110111101100","1001100011101001","1000101101001101","1001111111111010","1000111101100101","1000000001110010","1001110001110101","1001101010101101","1000000110010110","1010011001101001","1010011111010010","1000100011100111","1000111100111110","1000001111111011","1000011000100010","1000001110100101","1000010000001000","0000001110111100","0000100101101001","0000011010110011","0000011100101010","0000110010101100","0000011110110101","1000001111010011","1000000101011000","1000010001110111","1000001101110001","1000011011111000","1000001001001111","1000110100001000","1000011010010101","1010100011111011","1001010110100000","1000110010100001","1010000001011101","1010000111001000","1001101111011101","1000001100100111","0000001101101110","1000001100100100","1000010010101010","1000001101011010","1000010010100100","1000010000100001","1000101100011011","1000011111011001","1000001000001000","0000001100000000","0000001111101001","0000000111011010","0000001010001000","1000001010111110","1000010001101101","1000011011101101","1000000101101100","1000010100111110","1000011001111110","1001000010101001","1000011111110010","1011000101110010","1001000101001111","1000101110010100","1001101110010111","1000011111001011","1000010100001011","1000011000101001","0000001000000110","1000000001010111","0000000111110001","1000001011010100","1000011011110001","0000000011001100","1000011111001100","1000011001111110","1000100001011100","0000000011010011","0000010010111001","1000100111000110","1000010000000000","1000000011101101","1000011011110111","1000010000001010","1000010001110100","1000000001111011","1000100111010100","1000101011000111","1001010101010011","1011000100111101","1001001000001010","1000110001100011","1001010110101110","1010001110101010","1000001110011101","1000110010101001","0000001010110000","1000000100011000","1000000011000100","1000001011010111","1000001100110000","1000000011101011","1000000111101000","1000000110101000","1001001011011011","1000010011111001","1000010100011100","1000011111001111","1000010110011111","1000000100101011","1000000100110010","1000000100111101","1000001011010011","1000100010101011","1000011111101011","1001010100010000","1000010000000100","1010001000110011","1001001011100110","1001000000100100","1001100110100010","1000100110110000","1001001111101011","1000000101101010","0000011010010101","1000000111000001","0000011110001100","0000001100011110","0000001011010011","0000001000101101","0000001100110111","1000000101110111","1000101011011101","1000011100000010","0000000110110001","0000001101010000","0000110000010110","0000010111011100","0000000010001010","0000010000001000","0000001100101010","0000001000101010","1000100011000001","1001001000000110","1000011001110000","1001000110010011","1001010110110011","1000110010111111","1010100010001000","1000110001001011","1000010000111100","0000100001011110","0000010001111100","0000010101101101","0000010000100001","0000010110000000","0000011111101000","0000010010010011","0000001011001111","1000101010011000","1000011010001001","0000001100100110","0000010100101110","0000011001100000","0000100100000000","0000011010111110","0000010010001000","0000010001011110","0000010101100111","0000000111100100","0000011101100110","1000110010100010","1011100101011000","1011000010010010","1000111101100000","1000101101101000","1001111001110101","1000011101100001","1000011001010011","0001011010001111","0000001100011111","0000011010010011","0000100000010101","0000001001111110","0000000111001011","0000001000110101","1000010110101110","1000110011100100","1000001111111011","1000000011000110","0000010000001000","0000110001101000","0000100000101111","0000010110011010","0000011100011110","0000010000000001","0000001001011110","0000001001111110","1000111011110110","1001011001000000","1010001000101101","1000011001100110","1000110101000100","1000111000000111","1001011001001110","1000101101110101","0000100011000010","0000111111110011","1000000100111011","0000000100111110","0000010000001110","1000010111111011","0000001010001010","1000000110111110","1000100000101100","1000100000010000","1000011011110100","1000010101110000","0000001110111001","0000010001100110","0000010010000001","0000000101000100","1000001100110101","0000000000000000","0000010010101001","1000011001010110","1000111011100101","1010101011100100","1001010111001000","0000011011000010","1000010000101010","1000111000100101","1000000111001110","1001101111111110","1000010011101111","1000000101100110","1000000110010100","0000000110000110","1000000100100110","1000000111111011","1000010010011001","1000001010110000","1000001011010010","1000011001111010","1001000001100110","1000111101110010","1000000010001110","0000010101111010","0000011011110000","0000001000011011","1000000010001001","1000010010100110","1000001000111101","1000100100001110","1000010010010101","1010001110000110","1001010100100010","0000101100000011","1000111100010100","1000110000001100","1000111010010001","1001101101011110","1000101001011111","0000010101011111","1000100000111001","1000000100100010","0000001010101011","0000001001101001","1000011001000111","1000000111100101","1000001001111011","1000100010000111","1001000111011011","1000110010010010","1000011001111111","0000011001110000","0000010000001010","0000001100000010","1000010101101010","1000011110110100","1000100010111000","1000010100001111","1000010101010011","1001100000011000","1010110101101111","1000011001011110","1001000000101001","1000000100111100","1000111001111111","1000111101110111","1001000000001001","1000111001001000","1000010100101110","1000100101100111","0000010110001101","0000000010010011","1000011011011000","0000001111100110","1000000110001000","1000010101010100","1000100111111110","1000100111010011","0000001101101111","1000000110100100","0000001010000101","1000010101110001","1000011101010111","1000101011100111","1000011110001000","1001000111011101","1000110100000100","1001110000110101","1001010111100001","1001100000111111","1001011101011111","0000001100000110","1000101100011100","1000101110111111","1001110110111011","1001010000100100","1000110110000011","1000001001010111","1000010001101111","1000011110111011","1000010011101111","0000011010000001","1000000000110101","1001011101011110","1001010111101011","1000001100100101","1000000101010011","1000001001100010","0000000011100011","1000100000001110","1000101101110011","1000110011110010","1000111110110101","1000001111110111","1001010101100001","1010000110101101","1001010000100010","1001101001110001","1001010101110110","1000001010100010","1001001011010111","1010001001011101","1000110111011111","1001011010010011","1000100000010011","1000010111100101","0000000111000000","1000001111100000","1000110010010000","1000110011101110","1000110001001101","1000110001000011","1000110010110010","1000101010001111","1000110000110110","1000100000100010","1000110010011010","1000101111010010","1000001010000001","1000011100101111","1000101101011111","1000010100110000","1001011000000001","1001001111010110","1000110010111010","1001001100110001","1000110000001001","1000000101000101","1000111100000101","1000000111101111","1001111101111110","0000001010110110","1000001110111000","1000101111101000","1000101101101110","1000110110011100","1001100001000000","1001101111011110","1001111000110010","1010000011101100","1000111100010111","1001001011000110","1001001001101001","1000101110101010","1000101100101111","1000110011000110","1000001011100010","1000011111000000","1000110001000010","1001000001101011","1001000110111100","0000100001010101","0000101000111101","1001100111000010","1000000101010000","1000001000010111","1000111011100111","1001000100010010","1000110111001010","0000100000111001","0000010101000110","1000011111110111","1000100010110111","1000000101000101","1000100011011111","1000110100000101","1001011010010111","1001011000010100","1001010111001101","1001001111110100","1001001101100110","1000101011111101","1000111000010101","1001000100011000","1000110111101110","1000101011111010","1000011001100110","1001001010100011","1001010100111011","0000011011010100","1000010000100101","1000111101110101","0000000011111000","1000000100110101","1000000111010110","1010101111110101","0000010000010101","0000000111011001","1001001111111010","1000100110101111","1000010101010110","1000000100010000","1000000110001111","1000000110110011","1000100001011010","1000011101100000","1000111000101101","1000101010100011","1000111111000010","1000110000010000","1000110001100100","1000110011101010","1001001001111011","1000111111011000","1000110110000101","0000000011100011","1000001101011110","0000111011101010","1000001101001000","1001011100101110","1000000100010101","1000000011100001","1000000011010110","1001001000110001","1000011101010011","1000100010001001","1000101110111011","1000101011100111","1000001010110101","1000010100000111","1000100110100110","1000010110001100","1000100110011111","1000100011101010","1000110001110001","1000010000100001","1000110110111111","1000111010110011","1000100011101011","1000001010111001","1000010010011000","1000000110111000","1000010000011010","0000000111010111","0000000100111000","0000100101101000","1000110001100110","1001010010001001","1000000111100100","0000000011110000","0000000000101101","1001000000110001","1010100110011011","0000101000101001","1000000000011000","0000011010001000","0000010010111001","1000000111100111","1000010000110011","1000010011001101","1001000000000010","1000111001111110","1001001111001011","1001001100011101","1000011000011000","1000101000001100","1000010111101010","0000000000010001","1000000111000011","1000000101111010","1000000110011101","1000001100110011","0000110111101001","1000100011010010","1001000111000000","1000110101111011","0000000010000101","0000000001010111","0000000000010010","0000101101001101","1001110111011110","1000000100010101","0000011011011010","1000001011000000","0000000111001001","0000010010101010","0000000001001000","0000100000000110","1000010000111101","1000000101000001","0000000111011100","0000001110011100","1000001110011100","1000000000111100","0000011010000000","0000001011010111","0000001110000111","1000000011001001","0000010101011001","0000011001000010","1000111111000111","0000001110010011","1000000101110001","1000101100110001","1000000100010001","0000000011011010","0000000001010111","0000000011101001","0000110010010101","0000011110110101","0000100001111111","0000110011110110","0000101101101111","0000100011110111","0001000100101001","0000100101100110","0000100011000000","0000101101000110","0000011110011011","0001001100000000","0000010111000001","0000100101010100","0000100010100010","0000110010111101","0000101010011010","0000110101110010","0001010010010011","0000001010001011","0000110011000000","1000001101101100","1000101101011110","0000000000010011","1000000010111110","0000000110001110","1000000001000011","0000000101111111","1000000000011000","1001001011010100","1001011010011100","0000101001100001","0000000111111011","0000001100111011","0000001101000101","1000010110110110","1000001010111110","1000001001010010","1010111010000100","1000011101010010","1000001100000000","1001001101010110","1001001000100001","1000000100000101","1000011111110000","0000001100100100","0000010110010101","1000000001100111","1001001011111001","0000000011110100","1000000001111010","1000000001101101","1000000011100010");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
