library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_4 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_4;

architecture syn of ram_4 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"1000000000100111","0000000011101011","1000000010110010","0000000111010100","0000000010111010","1000000000100001","0000000010001111","0000000011011100","1000000011110110","0000000011101010","1000000100010110","1000000010111010","1000100100110111","1000101101010010","1000001010111001","1000000100100100","0000000010000101","1000000000111111","1000000001011011","0000000000110000","0000000100000010","1000000001101110","1000000010010001","1000000101010110","0000000111011001","1000000011010100","1000000000101001","1000000110011000","1000000001110101","1000000010111111","0000000101111100","0000000001100010","1000101001010000","1001001010100111","1001011010001010","1001110001101101","1001000001100000","1001110110101101","1001011110010000","1011010111011110","1011101111111000","1010000001000110","1000001100001011","1010000110100011","1010100011101100","1010110010000001","1011001011110010","1001101100101111","1001100111111000","1001011001101001","1001001010111011","1001010111111011","1000000010000111","0000000001100001","1000000111000100","1000000001111100","0000000000001111","0000000010010100","1000011111011010","1000110000101010","1001000010000111","1001000110110000","1001111100100010","1010100000110111","1001110011101011","1011000110001000","1011100000001101","1110010001100111","1100011001111001","1010011110000110","1001100001001011","1001101010000100","1001110101011000","1001000110111011","1011101001111101","1011100001111001","1010111011001000","1001010001100110","1001001110101010","1001011110000011","1010000100011001","1001000110010011","1000000000111111","1000000000110100","0000000000110110","0000000000111111","1000101011100110","1001001010100010","1000111101101101","1001000110010100","1001100101111001","1001011010001101","1010000011000010","1010100011110001","1001110010110001","1001110000110110","1100010100111000","1100110100101000","1011000111010000","1010101000111111","1010001111011110","1001100100100100","1001010001100110","1000110111000110","1000010000011100","1000010010001101","0000001010100111","1000011001101111","1000011000101011","1010000111110101","1000111001110001","1000000011000001","0000000111100101","1000000011101010","1000110001110110","1000111010011110","0000010000000000","0000001010101100","1000010000101000","1000001000110110","1000110111000000","1001001000011101","1001001111100011","1001011000001001","1001110101011110","1001011101110010","1001111101011011","1001101000111100","1001000110010111","1000100100101001","1000100111110101","0000001001010110","0000100000000000","0000010110100010","0000110110011110","0000010001010000","0001100111010000","0000011101100101","1000110100000100","1000110101011001","1000000011011111","0000000011110001","1001010000000011","1000111011000001","1000011100111110","0000100010110110","1000011011011011","1000100001110000","0000011000000000","1000000111100100","1000111101101111","1000110010101100","1000111000110001","1001101010000000","1000101010100000","1000100111001000","1000100111110111","1000001111110011","0000011111111101","1000100010100001","1000010011100110","1000110111100110","1000000001101011","0000010110111000","0000011111101001","1000010001011110","1001010001111110","1001011110101111","0000000000101000","1000000010100000","1001000110010011","1000110110000101","1000001001001101","1000000010110011","1001010111100001","1000100111110110","1000001100001100","1000010101001011","1000110101101110","1001000001000101","1001001111011101","1001101001010101","1001011101000001","1001110001111000","1001111010001000","1001010111101100","1000110101100110","1000111101001110","1000100001010011","1000010000000110","1000001110111001","0000100101000000","0000000110100001","1000100111101011","0000010000110100","1001111000100011","1000000000010000","1000110000100100","1001010111110111","1000100000010110","0000010011110010","0000110010101111","1000101010111110","1000100000100111","0000000001010000","1000010000011100","1000101000101110","1000011100110011","1001100010011000","1001011001010111","1001101100110111","1001110110111101","1001110010110100","1000110001110001","1000011100110110","1000100010101010","1000001110010011","1000010100001000","1000001110011011","0000000100110110","0000001110001111","1000100001111010","0000110001100111","1001111010010111","1000110111111111","1001000000010010","0000010011001100","1000010111001001","1000011010101111","1000011011110100","1000010010110000","1000010010100000","1000010111000111","1000100001000010","1000101110011001","1000100001101100","1001011011111001","1001011111100011","1001101000011110","1001101000011100","1001011110010000","1000110010100001","1000010010011010","1000110000011101","1000100001001001","0000001010110110","1000011101101101","1000010001011011","0000000101100010","0000000101100000","1000010011110101","1000111100110101","1000101011001010","1001100000110000","1000001101000010","1001110111110000","1001011011110111","1001010010101101","1000101001110101","1000010000010011","1000010001011001","1000101101001010","1000101110011110","1000101011111011","1000111100001010","1001000011000100","1010000010110111","1001110101011111","1000100101111000","1000011111011110","1000010110110111","1000110010110100","1000010010110101","1000001111101001","1000100000110011","1000000011010110","1001001111100000","1000101011100110","1001000000100000","1001100001100110","1000101000001100","1001011011100000","1001010101000110","1001101010001101","0000011010000100","1001000101010110","1000101100110011","1000010101010000","1000001110110101","1000001110100111","1000010110010111","1000011110111011","1000011010011010","1001011011110000","1010110000110001","1001010111100010","1000001101000111","1000000110101101","1000011100101110","1000010101110011","1000011000101001","1000010111111110","0000000010000010","1000111011011101","1000111111011101","1000101100000110","1001111101000110","1000110011000011","1000011011101110","1001001001111101","1001101011111100","1000011011110110","1001011001010100","1000100001101011","1000001100100110","1000100111000100","0000000100001011","0000001111110101","0000011101000011","0000000111110010","0000010001111011","1001110011010110","1010111000101110","1000110010011001","0000100100110011","0000010101111011","1000010100100111","1000011100110110","1000100000000011","1000110001110010","1000111000101011","1001100101100001","1010011100111101","1001011100111101","1001110111110000","1001000111010011","0000000010011100","1001000011110001","1001010011010101","1000011110101100","1001010111010101","1000100001000100","0000000111001111","0000010001111010","0000011111110101","0000001100100000","0000110001100001","0001000111101111","0001011100000111","1000011000100011","1001110110001111","1000010001000110","0000110111011000","0000011110100101","1000010011011101","0000000000000001","0000001010000100","0000001000101001","0000011100101011","1000101000100110","1000001100000011","1000101111111111","1001101101010101","1001010101001000","1000001001110010","1000011101100000","1001101001101100","1000100101011110","1000001101110100","0000000000111010","0000011111011011","0000010111011000","0000100111010100","0000100010110101","0000111000010001","0001000100001101","0000100110100101","1000100111110000","1000100110101111","1000000010100001","0000010111100111","0000010111111000","0000100101111110","1000000001010110","0000100011011111","0000101000110000","0000000111000101","1000011110100011","1001010000101110","1000110011100111","1000111111000101","1000110101000001","1000101101010001","1000001011011100","1001100001011010","1000001111101101","0000111110110001","0000100101101111","1000000010000110","0000100101100000","0000010100000100","0000010000011011","0000011001110011","0000011110101111","0000001111011001","1000100010101000","1000100101011010","1000010100101100","0000100111100110","0000111100101110","0000000101111100","0000011100101100","0000001001010111","1000000100101001","0000010101101011","1000010101100011","1000101111100110","1000010101010110","1010001001010010","1000111100001101","1000110011000111","0000001100110010","0001000000100001","0000001001100010","1000001001110001","1000010100011101","0000010011000001","0000100001100001","0000001000001010","0000011100100001","0000011101111100","0000010101011011","0000000001011000","1000100110000100","1000011100111111","0000010010001101","0001010100010110","0000101100101111","1000000101111011","0000010010000010","1000001010111000","1000001110011111","0000110001001011","1000010000101010","1001001110001110","1001000010100100","1000100010110000","1000000001101100","1000101001101011","1000001100000001","1000000000101000","1000101110110000","1000111110010000","1000010000000001","1000010011100010","0000100010010100","0000100001100100","0000001100010000","1000010011001011","1000001110000001","1000010100000100","1000010101010101","0000000101110001","0000101100001010","0000101010001111","0000100110011101","0000001111001110","0000001001001101","0000011100110010","0000010110110111","0000011001000000","1000000110100001","1000100110111010","1000111110011000","1001100111011011","1000010110000000","1000000010101111","1000001111100111","0000010111001101","1001011110111001","1000110110111011","1000100000101001","0000000101011110","0000010100011010","0000100101110000","0000001110111000","0000000101101110","1000011001010101","1000100010001111","0000001111101110","0000100011010101","0000011011001001","0000100000110101","0000011111000101","0000011100011111","1000011010001010","1000010100001010","0000000111110110","1000010100111101","1000001100111011","1001000000001010","1001011000011110","1001011000101000","1000110111100000","1000110110100111","1000001010001101","1000000000110001","1000100100101101","1000010111100011","1000010011001110","1000000001111010","0000000110011111","1000001110011000","1000001001011000","1000100100010100","1000101010101111","1000001100100110","0000001001011001","0000000111101111","0000011001010110","0000101001000100","1000101000110100","1000100011100111","1000011101000110","1000000111001011","0000011110101100","1000101001000110","1000001100010000","1001000110010101","1001011010110110","0000000010011110","0000101001001110","1000000101000001","1000111011100100","1000011000110100","0000010101111000","1000011100000110","0000001001111001","1000001111000100","1000011100011000","1000110000111001","1000111111010100","1000111011001011","1000110000011001","1001100011101010","1000100001011001","0000000101011101","1000001011100111","0000000001101011","1000100111011000","1000100011000100","1000110010000010","1000110010001111","0000011001001000","1001010011000001","1001011000110001","1001101001010100","1001111001110110","0000001110111100","1000011100010110","0000000100111110","1000111010010101","1000000010000110","1000000010011101","1001010011111111","1000101100010011","1001000000010001","1000110110010101","1001000011110000","1001100010110010","1001100111010101","1000111010110101","1001001000101010","1001000110011000","1000100100011010","1000001100011001","0000010011011111","0000001110101000","1000010000000001","1001000011110011","1001010011111001","1000011111111101","1001010111000000","1001011010101000","1000101101001001","1001010000011101","1001000001111111","1000101001111110","1000000101100001","1000000000101100","1000101100111101","1001000101110101","1001110101001111","1001000011010010","1010111001111111","1000110100011100","0000001110111001","1000011011101110","1000110001101111","1000111011111001","1001010000011000","1001010110101011","1001000011110011","1000100010011110","1000011011100100","0000000001110111","1000001011001100","1000000010111011","1000011110111000","0000001000110100","0000010111111001","1000000010010101","1000101011111110","1001000100000100","1000111001000100","1000000011111111","1000001011001000","1000001010100100","1000011010100011","1001001001000100","1001101111110100","1001000001110100","1000100011100010","1000110010001111","1000010100110111","1000101000001001","1000100000100001","1000110000111010","1001001011111110","1000111101111100","1001000111101100","1000110010101011","1000011101100100","0000000001100010","1000010110111010","0000110000000011","0000000011111011","0000001100001101","0000010011101111","0000001010011000","1000000011111001","1000110000000000","0000011010101001","1000000010100011","1000000100001001","1000000001100111","1000001111000111","1001001101101100","1010000010100010","1001011111110000","0000100111000000","0000100010111111","1000000001111100","0000001000000100","1000001110100011","1000100000010000","1000110101001011","1000110011110011","1000011101001011","1000010000111110","0000000001010011","0000001110100100","0000000100111010","0000101011111100","1000001011101110","0000011101010011","1000001011011001","1000111100011101","1001000010011010","0000011000101010","0000100000000011","1000000010101011","1000000011011010","0000000010001000","1000000101110100","1000101101001011","1001110010110100","0000010110111100","1000000100100100","1000000010110100","0000000100100011","0000100011001000","1000010111101011","1000001000100010","1000110100001100","1000101111001000","1000100110000110","1000010100000010","1000001100001001","1000001110001000","0000010010110010","0000011001101101","0000001110100000","0000001111110100","0000100011010010","0000110111101001","1000000110100000","0000101100001110","1000100001101000","1000000001100110","1000000000000010","0000000011001110","1000110111111111","1000000101100001","1001001101011110","1001110101011101","1000011000011101","1000111001101010","1000101110101001","1000010101100011","1000110110110100","1001000101010101","1010000101010101","1001001101010110","1001001010011110","1000100001101000","1001010000011101","1000111101000110","1000110000010011","1000111010010100","1000011110100010","1000010011111100","1000100001101110","0000001000001000","1000101001001111","1000111100110000","1000100111001100","0000000011010101","1000000011111101","0000000000010100","1000000010010001","1000100111001000","1001000101000010","1001000100100100","1010010001010000","1011101011111100","1001010000001010","1010100101100111","1010100000010000","1011010010100111","1010101111000101","1011110010111100","1101000010010111","1011110000011011","1011100011100010","1000111011110101","1010011010001000","1001011010111101","1001111101010111","1100000110101001","1010010110110010","1000101101110111","0000011110100110","1000001011110100","0000000011010101","1000000010011100","1000000001100101","0000000100001101","1000000010011010","0000000010011010","1000000011011110","1000001111001110","1000111011011111","1000111010000100","1001100111101110","1001100111111111","1001100011001000","1001011010001100","1001110101010010","1010010100100010","1010111100110101","1001100110000111","1001100011100010","1010010000001100","1010001100000011","1001000000100010","1001001111101011","1001000000011010","1000110100110001","1000001000100101","1000000010101100","0000000000111100","0000000101110001","0000000010100111");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
