library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_5 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_5;

architecture syn of ram_5 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"1000000010010111","0000000100011100","0000000011111010","1000000000000110","1000000100110011","1000000010110110","1000000011111010","1000000110010011","0000000010000110","0000000111001111","0000000000111111","0000000011101110","1000001101111111","1000010101000010","0000000010001110","0000000010111101","1000000111111111","1000000110000010","1000000110100001","0000000101101001","1000000111111100","1000000000000111","1000000010000010","1000000010001010","0000000011010111","0000000000011110","0000000101111001","0000000011100001","0000000000110000","0000000000011001","0000000000110010","0000000111001110","1000000001100100","1000000111110001","1000000100101101","1000001110110101","1000000110100010","1000010111000000","1000100011111000","1000101000011010","1000111101110111","1001001001100011","1010000110010101","1010011010111100","1010111000110010","1010100101101011","1001010000111010","1001010001101111","1001110011000011","1001001100110010","1000001110001000","1000000011010111","0000000000100101","1000000110000001","0000000110001010","1000000011011001","1000000001011110","0000000011100110","1000011010110100","1001001010101100","1001100111001111","1000110001100001","1000110101011010","1000110010101011","1001100111110011","1001110000001100","1001001111010100","1001001101111100","1001101100110110","1100001101011001","1011101100011000","1001101010010011","1000100010111111","0000000100010101","0000010101001011","0000001110010001","0000001111110101","1001101000000101","1000001110101100","1000000001110110","1001011100011101","1001000111011001","1000000100001101","0000000000010001","1000000000100100","0000000010111100","1000110100110110","0000011011100101","0000101101001111","1001000010111000","1001001000110100","1010101110001001","1010000101101101","1000111011010000","1000001101110101","1000011001101101","0000000110010100","1000000010100000","1000000100101111","0000000111000000","1000100100101110","1000001110111101","0000001010101110","0000011101110111","0000011000011001","0000011111100001","0000011100000110","1000001000000010","0000000101011111","1000010000110000","0000010000000000","0000000101000111","0000000010010110","1000101110000111","1001011011110110","0000010101111001","1010100100110111","1001001000111011","1000011101000101","1000001010110110","1001001111110001","1000111100100010","1000001100000001","0000001100100100","1000001001000111","1000111011001100","1000101100010100","1000001011011110","1000010111010101","1000001001011111","0000001110000000","1000001111001110","1000000111010100","0000011100110010","1000000000000111","0000001001010100","0000011100000100","0000011100111001","0001000110010001","1001001110101010","0000000000011001","0000000010100000","1001110110111001","0000011010010111","1010010010000111","1000101010001111","1000110010101001","1000101011000011","1000000011011110","1000000000010010","0000000111010011","0000010000110011","1000001010011100","1000001101010101","1000101110100000","1001000110101111","1000100010011010","1000001100101110","1000001101010111","1000001100000100","0000011111011111","0000001111010010","0000001010010111","0000010011000000","0000010001001110","0000110001110101","0000011000000011","1000111000110011","1000000010111001","1000101011111000","0000010110111101","1010101101001011","1000000000111011","1000001011100011","1000000100111010","1000011111000010","1000001100101100","1000000100110110","0000000010000110","0000000000101010","0000000011110110","1000011000100000","1000000101011110","1000110000010011","1000111011001011","1000101000111001","1000010100111110","0000010010110000","0000011011001010","0000001101101010","0000001000011000","0000011000101000","0000101000111011","0000100001101101","0000010000001011","1000000110011000","0000000000011010","1001101100110110","0000101000110000","1011101011111100","1010000011100001","1000010100011101","1000100100101101","1000000101011100","0000000111010101","1000001110100011","0000010011000111","0000011010011110","0000000010001011","1000011110110101","1000001111100001","1000111011100101","1000100000111111","1000100011110001","1000001001000000","1000001100111100","1000000011000111","0000000001011011","0000100110000010","0000001111000100","0000011001110110","0001011011010000","1000000000011000","1000000010101101","1000101011000000","1001010110011010","1010000101100110","1011110110001101","1001011000111000","1000000100011000","1000100110001010","1000000110001010","1000001110010110","1000000001111010","1000000001000001","0000011000111100","1000010010111000","1000101111100111","1000101100100111","1001001100000110","1000111010010011","1000101011100001","1000011111101110","0000000001110110","0000001000100101","0000000011001110","0000000001111110","0000101001010010","0001001101110010","0001000001010011","0000101001011000","1000001110001011","1000001000111100","1000111101111100","1001100010100000","1011101001101101","1001100101100000","1000010101111110","1000100110101011","1000010100101001","1000010101110111","1000011001110011","1000000100011010","0000101000100001","0000010011011100","1000100011000001","1001010111010110","1001111001010011","1001011110110100","1000111010110001","1000011001101001","1000001101101101","1000000011010100","0000011100111000","0000010100000101","0000100001110110","0001010110110010","0001100011101111","0000011110100000","1000010010000001","1000000101101101","1000111100011100","1001101010111001","1010100110111100","1000010000011110","1000010000010101","1000100110100111","0000000001100000","0000001001010111","0000010100100010","0000001111011000","0000001110110100","0000100111101011","0000000111000011","1000100111001110","1001001110000100","1001010000101000","1001011000011010","1001001001000111","1000110000110110","1000011101010001","0000000100001100","1000001011110010","0000010001010011","0010001110110001","0001000011001001","0001001101001010","1000111111010010","1000000110001110","1001011010010101","1010010000100001","1001011101001111","0000010001001010","1000011100000111","0000000011001010","1000000000101000","1000000001101101","1000010010101110","0000000011101110","0000011001011100","0000101000001011","0000101010110101","1000100010001001","1001001100100001","1001001001110000","1001000010001101","1000110100110101","1000111000011011","1001010111111100","1000111110111101","1000110111010101","0000011000010000","0010000100010101","0010010001111100","0001000010011110","1000101000011000","1000001011011010","1001001010001001","1010100000101110","0000011101111100","1000011010100110","1000100011110011","0000100000011011","0000000111001010","1000010010110101","1000010001000101","0000010000100000","0000011101010100","0000101010111111","0000010111101001","1000101100011100","1000111111011000","1001010010011101","1001010001100000","1001000000101101","1000111110111101","1001000110010011","1010011001110001","1010100011111111","1010100101000000","1011001101010010","1000110101001011","0001011111001101","1000111111101111","1000010001101001","1001000111100100","1001101011101110","0000011111101010","1000100100001011","0000100000101011","1000100010000001","1000000011011010","1000011111010011","0000000010101001","0000010111010111","0000100110110100","0000111000110111","0000000110011010","1000110100110100","1001011110011000","1001111110111010","1001001111111010","1000101101111001","1000100000011111","0000000000111100","1000101101100000","1000111100101101","1010001110101110","1011100011000110","1001111101001010","1000111001010001","1000110101000001","0000110000001011","1001000010101001","1001100000101001","1000010001001100","1000000010110011","1000010110110110","1000011101110100","1000011101010001","1000000100010110","0000001000011111","0000100001110011","0000010010111001","0000001011100100","1000011001101000","1000111000010011","1001010000110110","1001001010001101","1001000101010111","1000100110001111","1000101110001011","1000001100110010","0000000000100011","0000010100101000","0000111001001011","0000000101010011","1001001001101100","1001110010111110","1001001000000000","0000101110100000","1000100011011000","1001110110010111","1000110000010111","1000000110011110","1000110001011110","1000010110010111","1000110011111101","1000001010011000","0000000010001111","0000010010100010","0000010111110101","0000000101011011","1000101000111111","1001001011100111","1001011101011111","1001001001001001","1001000111000010","0000000101010100","1000000011110001","1000001101110101","0000100000110010","1000011001000010","0000011111111100","0001001111001110","0000010011111000","1010001000001100","1001011000000111","1000110000101110","1001001011010011","1010011000001000","0000000110100111","1000011011100101","0000000001111101","1000011101010000","1000111001100100","1000110100011011","1000110111110001","1000011111111011","1000010011100000","1000010011000101","1000110111100101","1001010001001101","1001000110011000","1001001101001110","1000111011000011","1000100000010100","1000000010101100","0000000010011100","0000001001010111","0000000100110100","0000010111000111","1000101110100100","0000001011011011","1010101111001101","1001001110000011","0000000101011001","1000110111011011","1010011000000110","0000100100100110","1000010001010100","0000011111100010","0000011010010110","1000100010100101","1000111010110010","1000110101010010","1001000101000100","1000110100010010","1001100111111001","1001110010010011","1001100110100011","1001000001010010","1000110000100101","1000001011101011","1000000100100001","1000001011111110","0000000100000010","0000000001010000","1000001100110011","0000010111110111","0000000010010101","1001000101011111","1010000000011110","1001010110011010","1001010011001001","1001010010101110","1010000001101111","0000011110000000","0000001001011010","0000100101100110","0000001111001110","0000001010101001","1000010111010110","1000011010000100","1000101001000011","1000001011011111","1000010100000001","1000100000001001","1000110001100011","1000111111100010","1000110010111011","1000001000101110","1000011000000101","1000010100111011","0000000100010010","1000001000111001","1000000111100010","0000000111111101","1000000000111000","1001010011000101","1010101001101011","1001010110111100","1000001011111100","1001011010010101","0000110000100101","0000011011101001","0000000100110010","0000000001100000","0000000111110111","1000010110100110","0000011001110001","0000000101100010","0000001011111110","0000001010000110","1000010101110000","1000101100011011","1000111000010010","1001000100110000","1001000010000101","1000011110101001","1000010100111110","1000010100101011","0000000000010011","1000000100110100","1000001000001001","0000100101100101","0000011100100001","0000100111111001","1010000011001000","1000111011100110","1000000000111110","1001100011101110","0000100111000000","1000001111001110","1000001011000111","0000010000000100","1000010001011111","1000000000100100","0000000110000111","0000001001100110","1000000101101101","0000011110010011","1000010100000101","1000100000001100","1000101000000000","1000110101111000","1000011010100101","1000010001000101","1000001010011000","1000000010110111","1000010101011100","1000001000100111","0000011011000111","0000010001011001","1000101001110101","0000000111000010","1001100100110010","0000110100100010","1000000111110010","1001101101000111","1010010110101010","0000100100010110","1000000000001100","0000000110110110","1000000000111111","0000010001111011","0000000100001110","0000000010011000","0000001101011111","0000010010001001","0000000111001000","1000000110011101","1000001001011010","1000010100010100","1000100110101001","1000001010110000","1000001101000111","1000010100110001","0000001101110100","0000010001001100","0000011010001101","1000001100011111","0000010000111110","0000100111011000","1000011000110100","1000011100111011","1000001100011011","1000011010101110","1011001001100001","0000100010001111","0000000110000111","1000011010011101","1000011001100000","1000010001001011","0000000011010111","1000001010011100","1000000011001100","1000001110011111","1000001001010111","1000000101110110","1000001010000111","1000100010000101","1000001100000011","1000001100110101","0000010001111010","0000001111010101","0000000101110001","1000000011000101","1000010001100010","0000110011000110","0000000111110010","1000000011011011","0000110001110110","1000101011010001","0000000011100001","0000000010111001","0000011111111101","0000111110111010","0000100000011001","1000001110011001","0000000001000101","1000010111100010","0000001011110101","1000000010011101","0000100011100001","1000001011000100","1000000110001011","1000001101101101","1000000001101000","1000001000010011","1000000000110011","1000011001001001","1000101001010010","1000000101001010","0000000011010001","1000001011111101","1000011101001100","0000110110001010","1000010110111010","1000100011100001","0000110010011010","1000000101111110","1000000100110001","1000000011111011","1010000100110110","0000010000001100","0000101000010000","1000001111110011","1000010000111001","1000001111111001","0000000110011110","0000011101010001","1000010001111100","0000000001001000","0000010011100100","0000100101101000","0000011011000111","0000000100011011","1000011010100011","0000000010000100","0000000110101010","1000010011000000","1000000101001011","1000011111110011","0000100110010101","0000010001001101","0000110001011011","1001101101000111","1000110100100111","0000000110110011","0000000011110101","0000000100101001","1000100010010010","0000101111000110","0000100001000100","0000000101110110","1000000001101101","1000010101111001","1000101110000100","0000101000000011","0000011010111001","0000000100111110","0000010111000101","0000101010101100","1000001110110000","0000101011100101","0000100000010001","0000110011010000","0000111000010111","0000011010001011","1000001101100110","0001001100011000","0001001111010010","0001010001001111","0001000001101011","1000001110010000","1000001101110001","0000000100000101","0000000000100011","0000000010100100","1000000100101011","1000011001110100","1001001001001101","1010011011101001","1010100110011111","1001010000111001","1001100010011101","1000111000010000","1000011110101111","0000011000011111","0000000100001010","1000100111000000","1000111101011100","0000010011100111","1000001101011101","1000101100101110","1000001111001111","1000000100111010","0000010011110111","0000111000111010","0001000011011010","1000110100001001","1000110100101101","1000000100100000","1000000101101111","1000000011001110","0000000001111111","0000000000001111","0000000010111001","0000000010100100","1000000110011101","1000000111101101","1000111001101011","1001010111111001","1001011011010111","1001010010110111","0000100001101000","0000100110011111","0000000010010101","1001000010110100","1010010111000110","1011111010011100","1010010111111100","1010010010110000","1001010011000111","1001010110010011","1001010101010000","1001010101010011","1000111101011111","1000110110111011","0000000101101000","1000000001011100","0000000010011000","0000000000101011");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
