library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_8 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_8;

architecture syn of ram_8 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"1000000001000111","1000000010001100","0000000000101001","1000000001001010","0000000001100101","1000000001110000","0000000100000001","0000000000000010","0000000001101101","0000000000000111","1000000010100011","1000000010001011","1000001000010000","1000011010111110","1000000101010000","1000000001011110","0000000011100100","0000000001001011","0000000001001100","1000000100110110","0000000111001101","0000000011100111","0000000010001100","0000000000100001","1000000010010101","1000000001001010","1000000110111011","0000000011100101","1000000011001000","0000000000101010","1000000001101010","0000000000110101","0000000000100000","0000000001001000","0000000010010100","1000001100110011","1000011101000011","1000011101110101","1000101100101000","1000110111101110","1000110111100101","1001000111000011","1001000000010101","1001100110111111","1001111110000100","1001110010010111","1001110101100101","1001010111001010","1001010000101111","1000110011010010","1000100000011111","1000001000100110","0000000111010010","0000000011000011","1000000001110010","1000000110100100","1000000000110111","0000000010111000","1000001011111101","1000010101000011","1000011010010001","1000010100011110","1000011111100111","1001000110001110","1001111000110100","1010110110001100","1011101100001110","1011101110100010","1101001000001110","1101010000000111","1110101001100101","1110011010100000","1110111010111011","1000110011001001","1000001100000110","1011010101100110","1100111101110000","1010001111100001","1001010010011001","1001011000010010","1001101010000110","1001001001100111","0000000100110001","1000000011010001","1000000000101011","1000000111001100","1000111001010000","1001001100110001","1000101101010101","1001111110101000","1010001010000111","1010111000101111","1000101011110111","1000100011011110","1000001100010010","1000011100101001","1000100111111000","1000100110110010","1000110011011111","1000101000110011","1000110101110010","0000000010111111","0000010010011101","1000111110011010","1000101111010011","0000000000111010","1000000010110110","0000011010100001","1000100010110111","0000000000001100","1000111011000001","0000000101001101","1000000000011100","1000000000010110","0000100010111100","1001011101111001","1001111100001000","1000110011110011","1001000100011100","1001001010101100","1000010000101101","0000011100001101","0000000111100001","0000000110001101","0000010111010010","0000001011001010","0000110011001110","0000000010011011","0000001010111100","0000001010000000","0000000111111100","1000010010001000","0000001110001101","0000001101001111","1000000100111101","1000011000110000","0000001010101101","0000101110010101","0000100111110010","1000001000111110","0000000011111101","0000000010100111","1001010101011110","1010010100011111","1001101001000110","1010001110100001","0000010101001100","1000000011011000","1000010101100101","1000000101011010","1000011000010010","0000010101101001","0000011100001001","0000001011101010","0000011110101110","1000001011000110","1000000011011010","0000001100100100","1000000001101110","1000001100000101","0000000110101100","0000000001001110","0000000010111001","1000100000101010","1000001011101101","0000001111111110","1000001001011010","1000011010111010","1000000011100100","1000010100110000","1010000010110000","1010111110100010","1000000101001111","1000011110111001","1000101000100010","1000000000001001","1000010000001011","1000001010011111","1000010010011010","0000000111100100","0000011001001011","1000000110101001","1000000111011110","0000001110100011","0000000010000001","1000000001001101","1000011000111111","0000000000100111","0000011010010101","1000000110101100","1000000100100001","0000010011100011","0000000000101000","0000100110100000","0000001100011111","1000100001111010","1000000011001100","1001011010101001","1010011000111111","1010000111001111","0000011111001111","1000010000100001","1000010011111100","1000000100011101","1000001101010101","1000000110010101","1000000001010000","1000001011001100","1000010011010100","1000010011001111","1000101110000100","0000010100000010","1000000111110000","1000100001111111","1000000000010101","0000000001100000","1000000011100100","0000000001100111","0000001010011001","0000000111110001","0000000011011111","1000010000110101","0000000010001101","1000100111001010","1000111011101101","1001110010110001","1010110011100000","1000000010110011","1000011001111011","0000000010111010","1000000000011100","0000000001100011","1000001000110000","0000000011100000","1000001010101111","1000000000101010","0000001111110100","0000001000100100","1000111111101000","1000100100100011","0000000110101100","1000011100101111","1000001101010011","0000001000101101","1000000001000110","1000000100010011","0000100101111000","0000001101110100","0000100000011000","0000010111010101","0000011101011011","0000101000100000","1000001110101011","1001011011101101","1001111001111001","1000110100100000","1000100100110100","0000010111111011","0000001111011110","0000000000111101","0000000011000100","1000000001111111","1000001010000001","0000001010000001","0000000111100101","1000001010110000","1001001100001100","1001010100011000","1000101000000000","1000011000100000","1000011110110000","0000000010010111","0000010011010011","0000010111101011","0000001001111001","0000000101010111","0000000011100111","0000001011111010","0000100100110101","1000101111110011","1000001100001010","1001101011101110","1010001011100001","1000111111100111","0000011101111100","1000010101111111","1000001010010010","0000000001011111","1000000100101100","1000001000100100","0000010110000101","0000001010100001","0000101111011001","1000000001100011","1000100111000010","1001001011111110","1001000101001011","1000110001100010","1000000100101000","0000001101000110","0000001000101010","0000000010000000","0000001110100000","0000011100110101","1000001101010101","1000100011010010","1000001111011110","1000001101101010","1000001001000011","1001101100101000","1010101100011111","1000011111000001","1000010001001010","1000010001011111","1000000010000000","0000010101010100","0000010010110000","0000001100111011","0000001110100101","0000010010100000","0000100101001110","0000101111001110","0000100011100100","1000011111111101","1000111001001100","1000101111100101","1000011001001110","1000010011001011","0000000110111010","1000000111101111","0000010111010101","1000010011101010","0000010100101001","1000100101100100","0001001010101001","1000001100011001","1000001110011111","1001000000010111","1001001100010111","1000001110011111","1000000110101001","0000001100010101","0000001001001110","1000001001110001","1000001100001111","1000001100110001","1000011000100111","1000010011100100","0000011101100101","0000101010000110","0000001001111001","1000010111111100","1000010111000001","1000001110001011","1000011001110110","0000001001000101","0000010010110100","0000100101011101","0000000011110110","0000100001100100","0000101010101011","1000010100000000","1000100111000110","1000011110100011","1000101010001111","1000110000011110","1001001110100100","1000101010010000","1000011011010011","1000100000111001","1000001111100010","1000001010100010","1000000001010111","1000001111100010","1000101111011100","0000000100100000","0000101001010110","0000101000010011","1000001100000010","0000000110001101","0000000100101000","1000101001001011","1000011010101100","1000000010000010","0000010011000101","1000000110111100","0000001111010111","0000001000100100","0000001100111001","0000001000110010","1000100100011011","0000001010100011","1000110010011101","1000111110111111","1001000100010000","1001000110111111","1001010011111010","1000100101101100","1000000110101101","1001010101111001","1000100011011111","1000111100101111","1000011000010010","0000101001101010","0000110100011001","0000011010011110","1000000110011100","1000010001000110","1000010100010111","1000010101111011","1000100100110010","0000000010011001","1000011110000011","1000001101110111","1000101010100110","1000111111110000","1000101110111100","0000101100011101","1000100001011111","1001000010111111","1000110100011110","1000011101111110","1001100111011001","1000011110011011","1001000100110101","1000111010001010","1001001000001111","1000110000111000","1000101110100011","1000010101100111","1000011011010011","1000000110010010","0000100001111011","0000011011110011","0000010011010011","1000010010011010","1000100110110010","1000100100000001","1000010101001110","1000010011110001","1000100110011111","1000100100100001","1000000001010001","1000011110011000","1000110100001000","0000000101100011","1001101110001011","1001000110001011","1000110010101111","1000111101001101","1001100110000010","0000000101011010","1001010110011101","1000110000001110","1000100001000100","1000011001001101","1000001111110011","1000011010110111","0000001110010101","1000000110000100","0000100101100011","0000000011001010","1000010111010010","1000010011010111","1000001010111111","1000011011000100","1000110001101100","1000111100111100","1000110110110101","1000101101101100","1000111010011001","1000011111110101","1000001011111000","1000101001101100","1010010011110110","1001000011011011","0000000101111010","1001011001111000","1000010110001111","1000001110100101","1000101101010001","1000111110111000","1000010011100111","1000001010011010","0000000101000100","0000001010111101","0000000111111101","0000011111010111","0000101110100110","0000000110110100","1000100011001011","1000110010011001","1000000101111010","1000110101011000","1001000011111110","1000101011110011","1000010000010011","1000000010011110","1000001101001101","0000010010101110","0000110110000110","1001000110101111","1001011111001000","1001110011011010","1000111001111010","1001000100010010","1000011100001110","1010100000110100","1000101000101100","1000010111111001","1000010001011001","1000010110001010","0000000011100010","0000000010000101","0000001010100110","0000010111100110","0000001101001111","1000001101010001","1000111110010111","1000101100110111","1000111101110110","1000111111111101","1000100100000110","1000001100111101","1000001011010101","1000010101111000","1000011000011110","1000011011100010","1000100011101000","1000010101101000","1001101110100110","1000111110001101","1000101010100100","1001100110001101","1010011111000010","1001010001111011","1000110101110000","0000011110001010","1000001111101010","1000011111101000","0000000111101100","1000000110001011","0000000011101101","1000100011001101","1000000101011011","1000101000111010","1001001001100111","1000101111010110","1000100110101111","1000011011101011","1000000101011111","1000001001101001","1000001100000100","1000011010001000","0000000110111001","0000011101001000","1000001100010011","1001100111000011","1010110001010110","1000111101110100","0000000001000110","1000111011000001","1010111101101110","1001000001001100","1000100111001001","1000010111000010","1000010010101011","1000000101011111","1000001011101111","1000010000100101","0000000001101001","1000111110001000","0000000000010100","1000010101111100","1001000110110000","1000010010011000","1000111010011010","1000010100010001","1000011010001010","1000001010101100","1000010000110100","0000001010100011","1000000001000110","0000000100110001","1000010011000111","1000110010000111","1001101000011101","1000110101101101","1000011101011100","1001010110101111","1010000001101001","1001010101001111","1000011100110000","1000100101011011","0000000101101010","0000000000001101","1000000100101110","1000000011110100","1000010100001111","1000100010101011","1000001000001100","1000001110011000","1000010110000000","1000011101101110","1000101010110000","1000010000110101","1000010011010011","1000000000010100","0000010001000110","0000000011001101","0000000111000110","1000001110110001","1001000001011101","1001001110101010","1001101110001011","1000100111100101","1000100000110101","1000100000100011","1001110111110001","0000001100001111","1000010011101100","0000000010000101","1000001001000000","1000000110100011","1000010100000010","1000011101011000","1000011101011111","1000001001001101","0000000000011111","0000000011010010","1000000000010000","1000011000010011","1000100101011011","1000010010101001","1000001100100000","1000011010010011","1000001100111100","1000001101100110","1000000010001101","1000010001001100","1000000101111101","1000000100001000","1001011110010000","1000101100000100","0000000011000001","0000000011011010","1001011110011010","0000001000111011","1000100001010001","1000101001001010","1000101010111101","1000011010111011","0000000101101000","1000101110010111","1000010011100010","0000000000000011","0000001000011001","0000011010101000","0000001011111000","1000000100010100","1000000101011001","1000001101111001","0000001010001101","1000000000111101","0000000010001000","0000000110010001","0000000011101010","0000011000011110","0000001011100111","1000100011000110","1001110001000100","0000000010001010","0000000001101100","1000000101110111","1000110101110001","1001101001111111","1010011001011110","1001001000000010","1000110000110001","1000100000110001","1000010011000110","1000010010111100","1000010101100110","0000011111011101","0000010111011011","0000001111000111","0000010011110111","0000010010100001","0000100001101001","1000101011000111","0000001010100000","0000101110100011","1000000100010000","1000100000111110","0000010101100001","1000110101011001","1000111011010000","1001011111011001","1001001010001001","1000000010000101","0000000011111100","0000000000110000","1000111000111101","1001010110010010","1010111010100001","1001000010000000","1000110110000101","1000111001110110","1000111100000010","1001010100001100","1000011101001101","1000011001010010","1001000001111010","1000101001001100","1000000111000100","0000010000011001","1000001001101100","0000000110000101","1000000111101001","0000011100101110","0000001011101001","1001100101110011","1010000111000011","1001000000010011","1001100111100101","1001000101001100","1000101111100100","0000000011111011","0000000111110000","1000000010001110","0000000001010110","1000101101010100","1010011101100010","1001101111010110","1010010001111011","1000111000000000","1000100011000001","1001110111101111","1001111010110110","1001100101011011","1001011100111001","1010000100000011","1010010101001001","1100110000011100","1101001010110000","1010011011100001","1001101000010011","1011001001111110","1010111000110111","1001100011001111","1001001011010001","1000010111011101","1000110010011001","1000010101001010","0000000101001100","0000000000110000","1000000001100011","1000000001011010","0000000000100111","0000000011001000","1000011101100001","1000100000100000","1001001110010011","1001111011001001","1010000010010110","1001111111000001","1001000100101100","1010001111100101","1010111011110000","1011011111110001","1011100001010101","1010010011010110","1010000111110001","1001111100011000","1001010100010100","1001010100101001","1001101111110010","1001100100000000","1001000100011101","1000110011000110","0000000011111001","1000000111101101","1000000011101010","1000000010111011");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
