library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_0 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_0;

architecture syn of ram_0 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"0000000101000010","0000000101000001","1000000010010110","0000000001000111","1000000001100101","1000000101011001","1000000001110001","1000000011000000","1000000010110001","1000000001111000","1000000110100111","0000000010000000","1000000100011001","1000000111101011","1000000001100100","1000000010100001","1000000011000010","1000000000010111","1000000101100011","1000000000010110","1000000010001000","1000000101100111","1000000110000011","0000000111101011","1000000111011110","0000000010101100","1000000011101000","0000000111011010","1000000110111100","1000000011110110","0000000010010001","0000000001100110","0000000010101111","1000000000101011","1000000100000101","1000000001101011","1000000111100101","1000100111001011","1000111000100000","0000101000101100","0000101101011110","0000101100010100","1010000111110111","1000101110011001","1000110011100100","1000101001100100","1001011000111001","1001000010101101","1000101001111101","1000101001010010","1000001010101100","1000000001110100","1000000111111000","1000000010100000","0000000011001010","0000000000000011","1000000011010110","0000000000111101","1000000111010010","0000110011001011","0000110111100110","1000111100111011","1000110110001000","0000000110100010","1001010010001011","1010011001000100","1010111010001000","1000110110111101","1000111111110011","1001101110011101","1011000100111101","1100001100111011","1010111111000010","1011101010111001","1100010100101001","1011011010000101","1011010100100000","1010110000100001","1001110010011001","1001011000101001","1000111100111010","1000010010011010","0000000001001010","0000000010001011","1000000010001101","0000000101110111","1000000000010110","0000100011111000","0000011001010111","1000101110001110","1001001001101100","1001001000111111","0000000111110010","1000110010010001","1000001100110111","1000000010011000","1000100110010111","1000001000110000","0000000001101111","1000011010011110","0000000111010011","0000001001110100","1000101010011101","1001000111011100","1000101101001100","1000001101111000","1001001100001001","1000011111111001","1000100111011000","0000010001110000","1000110110110100","0000000011011011","0000000110001011","0000000010110011","1000011110011111","1000001010110000","1000101011111000","1001011011111011","1001001000101001","1000100110000011","1000001111000011","0000011111111111","1000001110000000","0000001110011000","1000110011011000","1000001110010111","1000101001000101","1000010110011011","1000110011010101","1000010111100010","1000001110001011","0000101000100010","1000000101100110","1000101010000011","1000010101100011","0000101001100011","1000101011000010","1001000101011110","1001011010111110","1000000011111000","1000000001010101","1000000011010011","1001100010010111","1000100011000100","1001001011010011","1001100001010100","1000110010001110","1000110011110111","0000000010110100","1000000001101101","0000000000101101","1000001101101010","1000101101101110","1000000111101010","0000000000000101","1000010101100100","1000011001100001","1000000101100111","0000001111101101","0000010111100010","1000001011010101","1000100011111110","1000010000100101","1000010011100100","1000001101010001","1001111110001101","1010000111001111","1000111111101000","0000000011001100","1000000100010111","1001001001000111","1001010001011101","1000101100110001","1000101101001111","1000010010011101","1000010100101010","1000011110101011","1001001000011110","1000011010101010","1000010001100000","1000101011011111","1000000000000010","1000000000011101","1000011111011110","1000100000110100","1000010001100001","0000011100001111","0000001100110011","1000001111001011","0000010001100001","0000101000011011","1000000111000100","1001010001111111","1001101100000000","1001110100001010","1000011010011001","1000000101010000","1001001011010111","1000111110010101","1000101111001001","1000100111100100","0000011110101101","1000010100011110","1000100101100100","1000111111101000","1000000110111011","0000001000011101","1000000111101011","1000011010011111","1000010000111000","1000101010000010","1000010111101010","1000100001001001","0000001001000001","0000011011010101","0000011001011110","1000001001010001","1000011111010011","1000001010010111","0000010110101100","1000001000100000","1000100000100010","1001111000111110","0000010110101000","0000110001101111","1000111010111101","0000100011001100","0000111100000110","1001010011001001","1000101011001011","1000001000011000","1000110011011010","1000010001010101","0000000110110011","1000000100011101","1000011010110100","1000001010010101","1000010100010100","1000000100101001","1000000110111101","0000011110110111","0000001110101000","0000001011110000","1000000110011100","0000000010101100","0000001100010001","0000011001111010","0000101010011110","1000000100101000","1001101111100001","1010101101111110","1001011101000001","1000000011000110","1000101100001010","0001000000010111","0000011011110101","1001000001000100","1000000000010000","1000101000011001","1000111010110100","1000001110001010","0000001001011111","0000000010110101","1000100011111100","1000011010011100","0000000100110010","1000100100110111","1001000110110111","1000011011110100","0000000011000101","0000010100100001","0000011100011010","1000000110010100","1000011000110101","0000000010100100","0000011000001000","0000110111001100","1001111101111110","1010101110111011","1001001001011011","1000001010101101","1000011110000111","0000101100101010","0000101101110101","1000001000101011","0000111101011110","1000011000011110","1000011010001100","1000011000100010","1000001001100111","1000100111100001","1000000111110111","1000011000111011","1000011000011001","1000011110100100","1000111110100010","1000101001000010","0000000111100000","0000010000101011","0000000110010101","1000000110001111","1000000011111111","0000110010011111","0000101000011001","0000011110101000","1000111010011011","1010011100010000","1000010101101100","1000001010011010","0000110010001011","1001000001100010","1001110100100001","1001110000001001","1000111010111010","1000000101001101","1000001001011000","1000011100011011","1000010101111000","1000010010010101","1000001011110100","1000111011010010","1000011111101011","1001010100011000","1001111100011011","1001110000011001","1001000011101010","1000110001101100","0000001011101011","0000010011000010","0000100100010001","0000001101000001","0000100110001000","0000000111001111","1001010101100101","1010100101111110","1000011111010000","1000000111101000","0000101100110110","1000000010010011","1001011011001011","1001000101011101","0000001000101101","0000000111010110","1000010011100111","1000100101101111","0000001011100110","1000000101110111","1000000111110000","0000000111110001","1000100011000001","1010000101011110","1011000000010100","1010101001101111","1000111110100010","1000001101101111","0000001101010111","0000011001010011","0000001000011001","0000100110101001","0000011100011001","0000111110010101","1000001100110101","1001101011111001","1001000001001001","1000000111001001","0000110011111010","0000101011011100","1000111010010000","0000011101011100","0000000010100100","0000001000111100","0000001011010011","1000000010001100","0000000111011111","0000100001100111","0000000110010101","0000000001001010","1001101010100001","1010011100101111","1011010111010010","1010101001000011","1000011000010110","1000000101011011","1000010001000010","1000101001100011","1000000001011010","0000000000101010","0000111000001000","0000100001111110","1000000001001001","1001001111001110","1000110101011111","1000011111111111","1000001010111110","1000101011011011","1001100000100001","1000101110001111","0000011010100011","0000000111100110","0000100101111001","0000011000110000","0000100101110011","0000010111101110","0000010000000000","0000010011000100","1001010010011010","1011001111110000","1011011110101100","1010111000001111","1000010010101010","1000010011111011","1000010111001010","1000000000000111","0000100001110101","0000001111101101","0000101101010000","0000101111010101","0000000101000011","1001111100000110","1000110000100111","1000100100011001","1000000010011110","1001001001111100","1001110000010101","0000000001011001","0000001100010101","1000011110111000","0000011000101111","0000001111011000","0000101110010100","0000100110000100","0000001010101110","1000001110111001","1010010011001111","1011110001111100","1010110001000110","1001101111101011","1000111000001010","1000001111011100","1000001001000111","0000010110101110","0000001001000000","0000000100111000","0000101001111111","0000100100110100","0000100001100100","1001110001010011","1001001010111101","1000100000100111","1000001100010000","1001011101001111","1001010011011101","0000011000110001","0000011010010010","0000011010110010","0000000110111010","0000010100101100","0000100100101100","0000101001001101","0000011001001111","1001011011000000","1011110010110010","1011000101101001","1001011010101011","1001010011010000","1000011011111010","1000000110111011","1000000010110010","0000011010010100","0000000101000111","0000001010010000","0000000110110000","1000010001010000","1000011100111101","1001011100100110","0000100101000010","0000000011101011","1000011001000000","1001010111110000","1000100011101011","0000001110011001","0000011101010011","0000001111001001","0000001110011000","1000000111001011","0000101110001000","0001000001111111","0000000010000010","1001011001001111","1010101001111001","1010011011100100","1001100000010111","1000101010110101","1000001000011100","1000011000110101","1000000100110010","0000010001000101","1000001001000011","0000100000011101","0000001100001001","1000000100000111","1000100011011000","1001110111000110","0000110001111010","1000101111001100","1000010100001000","1001110011101001","1001010110010000","0000000001011111","1000000101100001","1000000010000000","0000010000101110","0000000011001000","0000100011110100","0000111010001001","0000000000111001","1001000010000111","1001110101101111","1001110111111000","1001001011100011","1000101111100010","1000011101111111","1000001000010010","1000000111100011","1000011110001111","1000001011011110","0000000110111011","0000010000111011","1000101111111111","1000010100011110","1001101011110000","1001000110001100","1000000010011101","0000101111101000","1000010101010101","1000110111110001","1000000100100001","1000100001011110","0000000111110101","0000000101110010","1000000000010111","0000000000011001","0000011000110110","0000010001100110","0000001011000101","1000111010010000","1001010101000101","1001001010001100","1000110011011101","1000010010101000","1000000100001101","1000010111100110","0000000001100111","0000001001001001","0000011011100001","0000000110000111","0000011000100010","1001100110100101","1010001110111001","1000100111001111","0000000100000111","0000101101101100","1000010000110111","1000010000010100","1000001110000010","0000100000010111","1000010101011001","0000000010011001","1000000011101111","0000001011101011","0000101001000000","0000101111010011","0000100101011011","1000001111010000","1000101101010111","1000011111111110","1000101010100001","1000011001000001","1000011101110111","1000010111010000","1000001100101010","0000011000011001","0000001001111100","1000111100011110","0000001000110010","1000111111010101","1000010001011010","1000001001011010","1000000001010010","1000110010110111","1000000101000011","1000000111110001","1000001000101110","0000010000010010","0000000111101001","0000000001111101","1000010001111000","0000000111101010","0000100111110100","0000110000000100","0000010100100001","1000010010101100","1000100010101000","1000010010101010","1000010110000000","1000101101111010","1000100111010100","1000110101011101","1000001111010110","1000000111010001","0000001100011101","1000101001011011","1000001101101010","1001000011000110","0000110001011011","0000101111100000","1000000010010010","1000000100010001","1001001110011111","1001010000011001","1001001001011010","1000001100000111","1000011101001111","1000100100111100","1000001001011110","0000000110000110","0000011011010011","0000001100011100","1000001011010111","0000010101110111","1000001010011001","1000010010110111","1000010001011010","1000001001011010","1000001100001101","1000001101010101","1000010010110001","0000000000100011","0000010111010011","0000000010011111","1001001010011010","0000010111100101","0000110100000100","0000101110100010","1000000111110101","1000000000001111","1000010000110011","1001111011001111","1001011010101100","1000100101111010","1000100010001110","1000000111111111","0000000000000110","0000100001000011","0001000001001101","0000101101010010","0000001011001111","0000000110100011","1000001100111100","1000010101000100","1000001010010100","0000001000000100","1000011111101001","1000111100110010","1001010001100000","1000110010011111","0000000111011100","1000101110001001","1001000001101101","1000000010101100","1000111010001010","0000000001111001","0000000001001111","1000000100010110","1000110000000111","1000110000011011","0000010000111110","1000011001110001","1000111100000101","1000101010111010","0000000110000010","0000101101011100","0000100000000010","0000000010001101","0000001101010101","0000001001011101","1000000010010011","0000000001000101","1000011110100101","1000001100011010","1000010100101100","1001011110001010","1010001100111011","1010000000101011","1000101011111011","1001000111001000","0000000110110001","1000000001010010","1000000001011111","0000000010000010","1000000110110111","0000000001101111","1000011100001011","1000001001110010","1000111000000100","1001110110111101","1001111000110101","1010000001001011","1010000010101011","1010101111100100","1011010001001100","1010011100100000","1011010001110100","1011011101111101","1011101000100000","1011000010100101","1010110010010100","1010111100011011","1011100100100001","1011101101100010","1010011000101001","1010000111000100","1001101011010011","1001001101001011","1000111111100110","0000000001111010","0000000001111101","0000000001010010","1000000010010101","1000000101101011","1000000001110011","0000000010011100","1000010100001001","1001010100011100","1001110000001100","1001011110010111","1010011000011111","1011100001110001","1011110010110101","1100001001001001","1100001111000110","1011001101101001","1010111110011111","1010101110011000","1010101010001100","1010011011101001","1010011100110110","1010011011111111","1001000011000110","1001000101011000","1000111100111110","1000101100010111","1000001111100110","1000001010011000","0000000010010011","1000000100001011","1000000001110011","0000000011000001","0000000011110011","1000000101010011","1000000001000111","1000011010100100","1000101001001100","1000110110111011","1000111101001011","1001001011111111","1001011010100111","1001001000100100","1001010010001010","1001001100110001","1010000010011001","1001100011111011","1001100110110010","1001001100101111","1000110010010010","1000010101110001","1000011111011100","1000110111011011","1000110011000100","1000101100011111","0000000000000001","0000000110101101","0000000010010111","0000000010010001");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
