library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_6 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(9 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_6;

architecture syn of ram_6 is

    type ram_type is array (0 to 783) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"0000000111111110","0000000011001010","1000000000111001","1000000011001011","0000000111111010","0000000001000101","0000000110001111","1000000100111011","1000000010101001","1000000010000000","0000000010110101","0000000011000111","0000100100111010","0000101010000101","1000101001111001","1000000111110000","1000000101011000","1000000011010110","0000000001011000","0000000000110100","0000000001001111","0000000000010101","1000000010001110","0000000001110111","0000000001000011","0000000011100011","1000000001001110","1000000011110111","0000000011010000","0000000001110000","1000000000111110","1000000001000111","0000100111000100","0001000011110011","0001010110110010","0001111010000110","0001000101001011","0001110110001010","0001011100100011","0001000110111101","0001100011101100","0001100001101011","1000011001001011","1000000011010110","1000101001000000","0001011101000010","0010001101101100","0010010110011011","0001100100110100","0001100101100001","0001000110111111","0001010100101100","1000000000111101","0000000110010001","0000000000110111","1000000011111000","1000000100001010","1000000001111111","0000100100111011","0000011010101011","0001000101101000","0000001011001110","0000011010111100","0001111010010110","0000111000100011","0000110000111110","0001011100110101","0001101001100100","0001010101110101","0000100000011001","0001001011101101","0000100111100000","0000110101101000","0001000010110001","0001001111100110","0001010101110101","0000100001010010","0010010001110110","0001010111010110","0000111000111100","0000010001110101","1000101000110010","1000000001001001","0000000001111101","1000000010111101","1000000000001000","1000110010010001","0000101000101111","1000101001111100","0000011011101010","0001001100011111","0000011111110010","1000001100101001","0000010010111010","0000111000001010","0000010001011011","0000010000010000","0000100101110111","0000001100100001","0000001100110101","0000000100111001","1000000100111100","0000011001110011","0000101001100100","0000010101110110","0000000011010011","0000110101000111","0000100111011010","0000011001000010","1000001011110011","0000010001111001","1000000010010000","1000000011011100","0000000011010111","1000110110111110","1000011111000000","1000011101100001","0000000100100001","1000100111001111","1000110011110011","1000011101000100","1000010100000001","0000001000100011","1000101000000000","1000101000100001","1000100101100101","1000100010110111","1000100101111111","1000010110101101","0000000000001011","1000000110100011","0000001001010110","0000100111001000","1000000011001001","0000100101011100","0000101010110111","1000010111111110","1000000001101000","1000010110110001","0000110101111100","0000000010101010","1000000000000000","0000101100010100","1001001100010011","1000100001010100","1001011110001000","1000101011101001","1000101011000110","1000011011011111","0000000011011101","0000010011110100","1001001011000011","1000101101110101","1001000111111100","1000100001101110","1000100000000011","1000101111110111","1000010000001000","1000000000110010","0000011001000010","0000010111000101","0000100110110100","1000000011010010","0000100101111011","0000101000001111","1000000101111101","0000100011110010","0000110010110000","0000000111100110","0000000000101001","0000010010010110","1000001110010100","1001001000001110","1000111110101100","1000010111001010","1000000011000001","1000100010100111","1000000100001000","1000100110010001","1000011111101001","1000100000101010","1000111000111101","1000101011110001","1000100111101010","1001000010010011","1000110110001011","1000110100100100","1000010101011010","1000000010101110","0000010111101110","0000010101100000","1000000101101101","0000100100100110","0000011110101101","1000100001011010","0000100001010101","0000000001001000","1000000010100011","1000110110010111","1000011111011111","1000111111111010","1001010010000100","1000110011000010","1000001010011000","1001000010001011","1000010001010100","1000011011011001","1000001011001001","1000011010010101","1000110100011111","1000100011010001","1000110100110111","1001010010010010","1000111111001111","1000110010110100","1000111110000100","1000010100011000","1000000110010011","0000000100010000","0000000000110011","0000110000001011","1000010101100000","0000000010111011","0000001100101101","1000101110011010","1000010011111101","1001000010111101","1010000100111010","1000101010011010","1001010110001010","1000101111111001","1000101110111100","1000110100111111","1000011110001101","1000100000100010","1000010100100001","1000100110100001","1000100101011100","1001000110000010","1001011101010010","1001011110000101","1001000110001011","1001100000001111","1001010110001111","1000101010001101","1000010010000110","1000001110101111","1000111010011101","1000110111111011","1000101000101111","1000100110111000","1001001001000111","0000000010001010","1000101011100010","1001011010000111","1000100010111010","0000011001111110","1001011000011100","1000101100100100","1000010001011000","1000110001000111","1000101010110111","1000110001001101","1000101111111001","1000101111101110","1001000010000001","1000110010110111","1001001010100100","1001010111101010","1001101111001101","1001011110001100","1001000001111101","1000011101111000","1000000000010100","1000011011010101","1000110100111000","1000100110001011","1001010101100000","1001011000110010","1001011011101110","1000000111100010","1000011001111010","1001000000110110","1000011011110101","1000101111000101","1000111101001101","1000111010111010","1000001111110110","1000100010010111","1000101111000101","1000010001100010","1000110001011001","1000100111010011","1000011010000000","1000111000111101","1001100011110110","1001010100001100","1001000101011110","1001001000110101","1001001010110110","1000011110101010","1000011011111110","1000111110110100","1000000001011101","1000001001101011","1001011100110001","1001100010011111","1000111000011111","1000000010101001","1000101101011001","1001010001101000","1001101001000111","1000101000110000","1000110111101111","1000110010011110","1000000000000101","1000101101011000","0000000000011111","1000010010011100","1000010111001010","0000001000101000","0000000100111110","1000111010101011","1001111100011101","1000111111010000","1001001110100101","1000111101001110","1000010110100100","1000000110011011","0000101010110001","1000000000110110","0000110101101000","1000001000111000","1001011101011001","1001110111110010","1000010111011011","0000000001100111","1000111000111000","1001010100100010","1001110101111111","1000100110101010","1000001101111000","1000000010111101","1000010110111000","1000010110101001","0000000111111010","1000000111010100","0000011101010000","0000010010011001","1000000011100111","1001001010001111","1001011000001111","1000101011100010","1000101101001111","1000011001000110","1000110000100101","1000000011101111","0000010000001100","0000100110100011","0001001010011111","0000100000001001","1000101100111110","1010010100011100","1000001001001100","1000010001001110","1000101101000000","1001100001011001","1010000111110011","1000101100000110","1000000111011101","0000000111001101","1000111100101111","1000010110110111","1000010011011111","0000100101001111","0000001111111101","0000001001011000","1000011001000010","1001000110111101","1000101101011011","1000010110000111","1000110000001101","1000100110010001","0000000100111100","0000001001000001","0000010001111100","0000110011110100","0001010100111110","0000110101011110","1000111000000101","1001111110100100","1000101010100010","1000001110001100","1000001101001010","1000001110001011","1010001010010111","1010001010010100","1000001010111110","0000000011010010","1000010100010010","1000000000101100","0000000110110110","0000110010110010","0000110001101001","1000000010000000","1000101010110100","1000101101110011","1000010100001011","1000010100110000","1001000000110010","1000011111000000","1000010011010011","0000001111011101","0000001100010111","0000101100100110","0000011101000001","0000011111001100","0000001000111011","1001010010111101","1001000101010111","1000001110010000","1000000000100010","1000011110111001","1010010100011100","1010100001011000","1000111011000110","0000000010011001","0000001100010000","1000000010000010","1000000010011000","0000010111101010","0000100011001010","0000001010011001","1000001010110000","1000001000011100","1000010101001000","1000100001101111","1000101010010110","1000001100110000","0000001010100000","0000001101010100","0000010100110001","0000010010110110","0000011011110000","0000011010101100","0000010110100111","1001000000001011","1001100000011000","1000000000001000","1000010001110000","1000110001011000","1001110101000101","1001000001010101","1000100001110011","1000001110101100","0000000110011010","0000010101110100","0000001101111010","0000100011101110","0001000110010011","1000011100110100","1000011011001000","1000001011110010","1000010110111110","1000101011100010","1000111111110011","1000000101111000","0000001100111100","1000001111110010","0000000000011101","0000011100111100","0000001101111100","0000011101100001","0000010001000101","1000110111111000","1001101010010001","1000000011010011","1000100100101000","1000110101101001","1001010100001010","1001100110001000","1000000011101111","1000010011111001","1000001101101111","0000011110001000","0000011000100111","0000110111110111","0001000111001110","1000011000001111","1000010011011100","1000010101111000","1000110001001000","1000111110000010","1000101001000110","1000011011101000","1000000101101001","0000000111010000","0000011101001100","0000011110000000","0000000001001000","1000000100001001","0000000011010101","1000110101000100","1010000010001010","1000001101010011","1000011011000111","1001010011000100","1000010101011100","1001000001000000","1001000111000111","1000001111110011","1000010000011111","1000000000010111","0000000001000011","0000100011100001","0000010100001101","0000101100001011","0000001100101110","1000011111000010","1000100110011001","1000010010111101","1000000110011000","0000000001111011","1000001111001100","1000001011001111","1000010101100001","0000000110010100","1000011001110110","1000010011101011","0000011000100011","1000011010010111","1001011000100111","1000001010111011","1000110100100001","1001010100100110","1001000011100100","1000100110111011","1001001001110001","1000100001010010","1000001111111011","1000101110000101","0000001000000011","0000011100100011","0001001100001110","0000100101101100","0000000110010110","0000000010110011","0000001001110110","1000001111100110","0000001011110100","0000001000000001","0000001111110011","0000001110000111","1000001110011111","0000010001010000","0000110110000011","1000011010000011","1001000111100001","1001010011010011","1001000001100111","1000000110110011","1000110001100100","1000110000101111","1011000000101011","1000110111110011","1000110110110001","1000101000001011","1000011010010010","1000101101011110","1000000011110010","0000100001100001","0000001110111000","0000011000111000","0000001010000100","0000100111011111","0000010010100011","1000000110001001","1000001000100110","0000001110110100","0000000100010010","0000100001101110","0000000001011111","1000010100000011","0000011101001111","1001001101110011","0000110010101001","1000011001111001","1000000110111100","1000001001100100","1000100010011000","1000110111100011","1001101101011101","1001101111110101","1001101001100110","1001010100010011","1000100110001110","1000010000001001","1000010110101101","0000000110111010","0000100010011110","0000111010101011","0000111111101100","0000011001100111","0000000011000010","1000001011010100","0000001010100011","0000100100010100","0000000111001110","0000011011000011","1000101010011111","0000010001110010","0000011000100010","1000101000010001","0000000110001001","1000011001100011","1000011101000101","1000000111100011","1000001111100010","1000001010011011","1001000010001100","1010110010100100","1011001011111011","1001010011100101","1000011101001011","1000110000111011","1000001011101101","0000010001111011","0000001010000011","0000001011011001","0000000001000101","1000010110100011","0000001010001101","1000010100001000","1000010001011000","1000010011011011","1000001000100001","0000000010111000","0000011111001000","1000100011110000","1000101101000010","1010000100011111","1000010111011110","0000101001111101","1000100101100000","1000000001100010","0000000111001001","1000000100001110","1000110100110010","1001000110100010","1001111001101100","1100101001111011","1010011010001001","1001010001010100","1000101110001110","1001001001100011","1001010001001010","1000111011100011","1000110000101101","1000101000011010","1000101011010010","1000110001101100","1000101000101000","1000000011110000","1000000010011000","0000001111000100","1000001010111110","1000001000100011","1011011100000100","1010000001111101","1001011101111111","1001011011001101","0000000101000101","0000000011001000","1000000001000010","0000000011000110","1000000100110111","1000011111100101","1001001110000111","1001111101011000","1011011110110100","1100010001111110","1101011001111111","1110011000011001","1011110000010011","1010110010100101","1010100110111100","1010010000101000","1001011100000011","1000100110111111","1001000001111101","1001011011000001","1010001001011011","1001110100101001","1100001110111010","1011010011010100","1001100111000001","1001001010011010","1000011010010110","1000001000111111","1000000000011011","0000000011000011","0000000000000000","0000000011001110","1000000100101001","1000011011100101","1000101000100010","1001001001011100","1001011111010000","1010011011110111","1010110010000010","1100101001001100","1001000111100011","1000010110000000","1011110011101011","1011100111100011","1011110101011110","1011110110011010","1100110100000001","1011111101011001","1010101001111011","1001110111111000","1001011011111000","1001000111010010","1000111010100000","1000100010111001","1000000101001110","1000000111000110","0000000000110010","0000000000101110","1000000001101011","1000000100110000","1000000001100000","1000000010111110","1000001110000011","1000001111101001","1000010110101011","1000101111010010","1001000101100111","1001100110100001","1010001111011001","1010101100100000","1001100010101111","1001101110100101","1011100000001110","1011011110000110","1010110010110110","1010001000001001","1001011010100010","1001001100010110","1001000011100110","1000100101011100","1000101000000101","1000010110110000","0000000000000010","1000000000101000","1000000000110110","0000000000101111","1000000011111101","1000000011010000","0000000010110110","1000000100101000","1000000110001011","1000001100111111","1000000000011110","1000000110001010","1000000000001011","1000010110111110","1000001101001000","1000011001101100","1000010111000100","1000100111110100","1000010001101110","1000010000000000","1000010100001011","1000010010111110","1000010001101110","1000001010011100","1000001100111101","1000010000000101","0000000000100110","1000000100000001","0000000001000111","0000000010110000","0000000010001110");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));
end syn;
